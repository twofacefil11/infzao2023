<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.698,-1.21657,47.8846,-46.8322</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>29,-11</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>29,-16</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>36.5,-14</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,-15</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>22.5,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>42,-14</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>16,-10</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>16,-12</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>45,-14</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-10,26,-10</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>20 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>20,-15,20,-10</points>
<intersection>-15 10</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-15,20.5,-15</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>20 9</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-17,19,-12</points>
<intersection>-17 3</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-12,26,-12</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>19 0</intersection>
<intersection>26 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19,-17,20.5,-17</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>26,-12,26,-12</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-13,32.5,-11</points>
<intersection>-13 1</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-13,33.5,-13</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,-11,32.5,-11</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-15,26,-15</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-17,26,-17</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-14,40,-14</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-16,32.5,-15</points>
<intersection>-16 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-16,32.5,-16</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-15,33.5,-15</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-14,44,-14</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 1>
<page 2>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 2>
<page 3>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 3>
<page 4>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 4>
<page 5>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 5>
<page 6>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 6>
<page 7>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 7>
<page 8>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 8>
<page 9>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 9></circuit>