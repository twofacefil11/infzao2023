<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport>
<gate>
<ID>1</ID>
<type>AA_REGISTER4</type>
<position>23,-23</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>7 </output>
<output>
<ID>OUT_2</ID>9 </output>
<output>
<ID>OUT_3</ID>10 </output>
<input>
<ID>clear</ID>6 </input>
<input>
<ID>clock</ID>5 </input>
<input>
<ID>count_enable</ID>11 </input>
<input>
<ID>count_up</ID>13 </input>
<input>
<ID>load</ID>12 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>2</ID>
<type>DD_KEYPAD_HEX</type>
<position>11.5,-22.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 10</lparam></gate>
<gate>
<ID>3</ID>
<type>CC_PULSE</type>
<position>19,-29.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>27,-29.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>33.5,-23</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>9 </input>
<input>
<ID>IN_3</ID>10 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>19,-12</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>23,-15</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>28,-15.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-21,17.5,-19.5</points>
<intersection>-21 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-19.5,17.5,-19.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-21,19,-21</points>
<connection>
<GID>1</GID>
<name>IN_3</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-21.5,19,-21.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-22,19,-21.5</points>
<connection>
<GID>1</GID>
<name>IN_2</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16.5,-23.5,19,-23.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-23.5,19,-23</points>
<connection>
<GID>1</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-25.5,17.5,-24</points>
<intersection>-25.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-24,19,-24</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-25.5,17.5,-25.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-29.5,22,-27</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-29.5,22,-29.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-29.5,24,-27</points>
<connection>
<GID>1</GID>
<name>clear</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-29.5,25,-29.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-23,30.5,-23</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-24,30.5,-24</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-22,30.5,-22</points>
<connection>
<GID>5</GID>
<name>IN_2</name></connection>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-21,30.5,-21</points>
<connection>
<GID>5</GID>
<name>IN_3</name></connection>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>23,-18,23,-17</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1</GID>
<name>count_enable</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-18,21,-12</points>
<intersection>-18 4</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-12,23,-12</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-13,23,-12</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21,-18,22,-18</points>
<connection>
<GID>1</GID>
<name>load</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-15.5,26,-15.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>24 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,-18,24,-15.5</points>
<connection>
<GID>1</GID>
<name>count_up</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 1>
<page 2>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 2>
<page 3>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 3>
<page 4>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 4>
<page 5>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 5>
<page 6>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 6>
<page 7>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 7>
<page 8>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 8>
<page 9>
<PageViewport>-0.0479392,0,44.2479,-46.2</PageViewport></page 9></circuit>