<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-15.6427,54.322,43.6166,-27.1308</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>14.5,28.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>9,3</position>
<input>
<ID>N_in3</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>20.5,19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_FULLADDER_4BIT</type>
<position>13.5,10</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>9 </input>
<input>
<ID>IN_B_0</ID>13 </input>
<input>
<ID>IN_B_1</ID>12 </input>
<input>
<ID>IN_B_2</ID>11 </input>
<input>
<ID>IN_B_3</ID>10 </input>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>5 </output>
<output>
<ID>OUT_2</ID>3 </output>
<output>
<ID>OUT_3</ID>2 </output>
<input>
<ID>carry_in</ID>18 </input>
<output>
<ID>overflow</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>16.5,28.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>18.5,28.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>20.5,28.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>33.5,33</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>-1.5,28.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>0.5,28.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>2.5,28.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>4.5,28.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>12,3</position>
<input>
<ID>N_in3</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>18,3</position>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>15,3</position>
<input>
<ID>N_in3</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AI_XOR2</type>
<position>25.5,19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>15.5,19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AI_XOR2</type>
<position>30.5,19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>3,6.5</position>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,4,9,6</points>
<connection>
<GID>4</GID>
<name>N_in3</name></connection>
<intersection>6 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,6,12,6</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,4,12,5</points>
<connection>
<GID>17</GID>
<name>N_in3</name></connection>
<intersection>5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13,5,13,6</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12,5,13,5</points>
<intersection>12 0</intersection>
<intersection>13 1</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,4,18,6</points>
<connection>
<GID>18</GID>
<name>N_in3</name></connection>
<intersection>6 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>15,6,18,6</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,4,15,5</points>
<connection>
<GID>19</GID>
<name>N_in3</name></connection>
<intersection>5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>14,5,14,6</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14,5,15,5</points>
<intersection>14 1</intersection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,14,11.5,17</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>17 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>4.5,17,4.5,26.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>17 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,17,11.5,17</points>
<intersection>4.5 1</intersection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,14,10.5,16</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2.5,16,2.5,26.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,16,10.5,16</points>
<intersection>2.5 1</intersection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,14,9.5,15</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>0.5,15,0.5,26.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0.5,15,9.5,15</points>
<intersection>0.5 1</intersection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-1.5,14,-1.5,26.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,14,8.5,14</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>-1.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,14,15.5,16.5</points>
<connection>
<GID>8</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,14,16.5,16</points>
<connection>
<GID>8</GID>
<name>IN_B_2</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16.5,16,20.5,16</points>
<intersection>16.5 0</intersection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,16,20.5,16.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>16 2</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,14,17.5,15</points>
<connection>
<GID>8</GID>
<name>IN_B_1</name></connection>
<intersection>15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,15,25.5,16.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17.5,15,25.5,15</points>
<intersection>17.5 0</intersection>
<intersection>25.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>30.5,14,30.5,16.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18.5,14,30.5,14</points>
<connection>
<GID>8</GID>
<name>IN_B_0</name></connection>
<intersection>30.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,22.5,14.5,26.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,22.5,19.5,23</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17.5,23,17.5,26.5</points>
<intersection>23 2</intersection>
<intersection>26.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17.5,23,19.5,23</points>
<intersection>17.5 1</intersection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16.5,26.5,17.5,26.5</points>
<intersection>16.5 4</intersection>
<intersection>17.5 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16.5,26.5,16.5,26.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>26.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,22.5,24.5,24</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>18.5,24,18.5,26.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18.5,24,24.5,24</points>
<intersection>18.5 1</intersection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,22.5,29.5,24.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>24.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20.5,24.5,20.5,26.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20.5,24.5,29.5,24.5</points>
<intersection>20.5 1</intersection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,25,33.5,31</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>25 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>16.5,22.5,16.5,25</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>16.5,25,33.5,25</points>
<intersection>16.5 1</intersection>
<intersection>21.5 9</intersection>
<intersection>26.5 4</intersection>
<intersection>31.5 5</intersection>
<intersection>33 3</intersection>
<intersection>33.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,11,33,25</points>
<intersection>11 7</intersection>
<intersection>25 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>26.5,22.5,26.5,25</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>25 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>31.5,22.5,31.5,25</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>21.5,11,33,11</points>
<connection>
<GID>8</GID>
<name>carry_in</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>21.5,22.5,21.5,25</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>25 2</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,7.5,3,9</points>
<connection>
<GID>23</GID>
<name>N_in3</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,9,5.5,9</points>
<connection>
<GID>8</GID>
<name>overflow</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 1>
<page 2>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 2>
<page 3>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 3>
<page 4>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 4>
<page 5>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 5>
<page 6>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 6>
<page 7>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 7>
<page 8>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 8>
<page 9>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 9></circuit>