<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>14.698,-1.21657,47.8846,-46.8322</PageViewport>
<gate>
<ID>10</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,-16</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,-19</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>16,-14</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>16,-21</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>44,-17.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>32,-15</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>32,-20</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>39,-17.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>31.5,-29.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>35.5,-29.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-28.5,23.5,-14</points>
<intersection>-28.5 12</intersection>
<intersection>-19 10</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-14,29,-14</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>23.5,-19,24,-19</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>23.5,-28.5,28.5,-28.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-21,22.5,-16</points>
<intersection>-21 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-21,29,-21</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>20 9</intersection>
<intersection>22.5 0</intersection>
<intersection>29 11</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-16,24,-16</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>20,-30.5,20,-21</points>
<intersection>-30.5 10</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-30.5,28.5,-30.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>20 9</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>29,-21,29,-21</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-21 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>42,-17.5,43,-17.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-16.5,35,-15</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-16.5,36,-16.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-20,35,-18.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-18.5,36,-18.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-16,29,-16</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-19,29,-19</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-29.5,34.5,-29.5</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<connection>
<GID>26</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 1>
<page 2>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 2>
<page 3>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 3>
<page 4>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 4>
<page 5>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 5>
<page 6>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 6>
<page 7>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 7>
<page 8>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 8>
<page 9>
<PageViewport>0,0,77.7,-106.8</PageViewport></page 9></circuit>