<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>7.10543e-015,-18.5625,139.4,-88.7625</PageViewport>
<gate>
<ID>2</ID>
<type>AA_RAM_4x4</type>
<position>70,-34.5</position>
<input>
<ID>ADDRESS_0</ID>4 </input>
<input>
<ID>ADDRESS_1</ID>3 </input>
<input>
<ID>ADDRESS_2</ID>2 </input>
<input>
<ID>ADDRESS_3</ID>1 </input>
<input>
<ID>DATA_IN_0</ID>10 </input>
<input>
<ID>DATA_IN_1</ID>9 </input>
<input>
<ID>DATA_IN_2</ID>8 </input>
<input>
<ID>DATA_IN_3</ID>11 </input>
<output>
<ID>DATA_OUT_0</ID>10 </output>
<output>
<ID>DATA_OUT_1</ID>9 </output>
<output>
<ID>DATA_OUT_2</ID>8 </output>
<output>
<ID>DATA_OUT_3</ID>11 </output>
<input>
<ID>ENABLE_0</ID>7 </input>
<input>
<ID>write_clock</ID>5 </input>
<input>
<ID>write_enable</ID>6 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:8 11</lparam>
<lparam>Address:9 15</lparam>
<lparam>Address:15 1</lparam></gate>
<gate>
<ID>10</ID>
<type>DD_KEYPAD_HEX</type>
<position>57.5,-34.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>14</ID>
<type>CC_PULSE</type>
<position>73,-29</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>80,-36</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>86,-35</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>70,-46</position>
<input>
<ID>ENABLE_0</ID>6 </input>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>15 </input>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>8 </output>
<output>
<ID>OUT_3</ID>11 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>73,-51</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_TOGGLE</type>
<position>71,-51</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>69,-51</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>67,-51</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>55,-51</position>
<input>
<ID>N_in3</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>57.5,-51</position>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>60,-51</position>
<input>
<ID>N_in3</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>62.5,-51</position>
<input>
<ID>N_in3</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-33,63.5,-31.5</points>
<intersection>-33 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-33,65,-33</points>
<connection>
<GID>2</GID>
<name>ADDRESS_3</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-31.5,63.5,-31.5</points>
<connection>
<GID>10</GID>
<name>OUT_3</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-34,63.5,-33.5</points>
<intersection>-34 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-34,65,-34</points>
<connection>
<GID>2</GID>
<name>ADDRESS_2</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-33.5,63.5,-33.5</points>
<connection>
<GID>10</GID>
<name>OUT_2</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-35.5,63.5,-35</points>
<intersection>-35.5 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-35,65,-35</points>
<connection>
<GID>2</GID>
<name>ADDRESS_1</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-35.5,63.5,-35.5</points>
<connection>
<GID>10</GID>
<name>OUT_1</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-37.5,63.5,-36</points>
<intersection>-37.5 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-36,65,-36</points>
<connection>
<GID>2</GID>
<name>ADDRESS_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-37.5,63.5,-37.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-33,76,-29</points>
<intersection>-33 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-33,76,-33</points>
<connection>
<GID>2</GID>
<name>write_clock</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-29,76,-29</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-34,83,-34</points>
<connection>
<GID>2</GID>
<name>write_enable</name></connection>
<intersection>83 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>83,-44.5,83,-34</points>
<intersection>-44.5 15</intersection>
<intersection>-36 13</intersection>
<intersection>-35 12</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>83,-35,84,-35</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>83 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>82,-36,83,-36</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>83 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>67,-44.5,83,-44.5</points>
<intersection>67 16</intersection>
<intersection>83 10</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>67,-46,67,-44.5</points>
<connection>
<GID>24</GID>
<name>ENABLE_0</name></connection>
<intersection>-44.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-36,76.5,-35</points>
<intersection>-36 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-35,76.5,-35</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-36,78,-36</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-44,69.5,-39.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>-42 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>57.5,-42,69.5,-42</points>
<intersection>57.5 9</intersection>
<intersection>69.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>57.5,-50,57.5,-42</points>
<connection>
<GID>33</GID>
<name>N_in3</name></connection>
<intersection>-42 8</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-44,70.5,-39.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>-42.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>60,-42.5,70.5,-42.5</points>
<intersection>60 9</intersection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>60,-50,60,-42.5</points>
<connection>
<GID>34</GID>
<name>N_in3</name></connection>
<intersection>-42.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-44,71.5,-39.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-43 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>62.5,-43,71.5,-43</points>
<intersection>62.5 9</intersection>
<intersection>71.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>62.5,-50,62.5,-43</points>
<connection>
<GID>35</GID>
<name>N_in3</name></connection>
<intersection>-43 8</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-44,68.5,-39.5</points>
<connection>
<GID>2</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>-41.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>55,-41.5,68.5,-41.5</points>
<intersection>55 9</intersection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>55,-50,55,-41.5</points>
<connection>
<GID>31</GID>
<name>N_in3</name></connection>
<intersection>-41.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-49,73,-48</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-48,73,-48</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-49,71,-48</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-48 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-48,71,-48</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-49,69,-48</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-48,69.5,-48</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-49,67,-48</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-48,68.5,-48</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>17.425,-8.775,121.975,-61.425</PageViewport>
<gate>
<ID>36</ID>
<type>AA_RAM_4x4</type>
<position>68.5,-27.5</position>
<input>
<ID>ADDRESS_0</ID>20 </input>
<input>
<ID>ADDRESS_1</ID>19 </input>
<input>
<ID>ADDRESS_2</ID>18 </input>
<input>
<ID>ADDRESS_3</ID>17 </input>
<input>
<ID>DATA_IN_0</ID>26 </input>
<input>
<ID>DATA_IN_1</ID>25 </input>
<input>
<ID>DATA_IN_2</ID>24 </input>
<input>
<ID>DATA_IN_3</ID>27 </input>
<output>
<ID>DATA_OUT_0</ID>26 </output>
<output>
<ID>DATA_OUT_1</ID>25 </output>
<output>
<ID>DATA_OUT_2</ID>24 </output>
<output>
<ID>DATA_OUT_3</ID>27 </output>
<input>
<ID>ENABLE_0</ID>23 </input>
<input>
<ID>write_clock</ID>21 </input>
<input>
<ID>write_enable</ID>22 </input>
<gparam>angle 0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:5 5</lparam>
<lparam>Address:6 6</lparam>
<lparam>Address:8 8</lparam>
<lparam>Address:9 9</lparam>
<lparam>Address:11 10</lparam></gate>
<gate>
<ID>37</ID>
<type>DD_KEYPAD_HEX</type>
<position>56,-27.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<output>
<ID>OUT_1</ID>19 </output>
<output>
<ID>OUT_2</ID>18 </output>
<output>
<ID>OUT_3</ID>17 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>38</ID>
<type>CC_PULSE</type>
<position>71.5,-22</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AE_SMALL_INVERTER</type>
<position>78.5,-29</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>84.5,-28</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>68.5,-39</position>
<input>
<ID>ENABLE_0</ID>22 </input>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<input>
<ID>IN_2</ID>34 </input>
<input>
<ID>IN_3</ID>35 </input>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>25 </output>
<output>
<ID>OUT_2</ID>24 </output>
<output>
<ID>OUT_3</ID>27 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>53.5,-44</position>
<input>
<ID>N_in2</ID>40 </input>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>56,-44</position>
<input>
<ID>N_in2</ID>42 </input>
<input>
<ID>N_in3</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>58.5,-44</position>
<input>
<ID>N_in2</ID>43 </input>
<input>
<ID>N_in3</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>61,-44</position>
<input>
<ID>N_in2</ID>41 </input>
<input>
<ID>N_in3</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>DD_KEYPAD_HEX</type>
<position>68.5,-51.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<output>
<ID>OUT_1</ID>33 </output>
<output>
<ID>OUT_2</ID>34 </output>
<output>
<ID>OUT_3</ID>35 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>55</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>58.5,-52</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>40 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 8</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-26,62,-24.5</points>
<intersection>-26 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-26,63.5,-26</points>
<connection>
<GID>36</GID>
<name>ADDRESS_3</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-24.5,62,-24.5</points>
<connection>
<GID>37</GID>
<name>OUT_3</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-27,62,-26.5</points>
<intersection>-27 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-27,63.5,-27</points>
<connection>
<GID>36</GID>
<name>ADDRESS_2</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-26.5,62,-26.5</points>
<connection>
<GID>37</GID>
<name>OUT_2</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-28.5,62,-28</points>
<intersection>-28.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-28,63.5,-28</points>
<connection>
<GID>36</GID>
<name>ADDRESS_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-28.5,62,-28.5</points>
<connection>
<GID>37</GID>
<name>OUT_1</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-30.5,62,-29</points>
<intersection>-30.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-29,63.5,-29</points>
<connection>
<GID>36</GID>
<name>ADDRESS_0</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-30.5,62,-30.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-26,74.5,-22</points>
<intersection>-26 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-26,74.5,-26</points>
<connection>
<GID>36</GID>
<name>write_clock</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-22,74.5,-22</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-27,81.5,-27</points>
<connection>
<GID>36</GID>
<name>write_enable</name></connection>
<intersection>81.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>81.5,-37.5,81.5,-27</points>
<intersection>-37.5 15</intersection>
<intersection>-29 13</intersection>
<intersection>-28 12</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>81.5,-28,82.5,-28</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>81.5 10</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>80.5,-29,81.5,-29</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>81.5 10</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>65.5,-37.5,81.5,-37.5</points>
<intersection>65.5 16</intersection>
<intersection>81.5 10</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>65.5,-39,65.5,-37.5</points>
<connection>
<GID>41</GID>
<name>ENABLE_0</name></connection>
<intersection>-37.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-29,75,-28</points>
<intersection>-29 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-28,75,-28</points>
<connection>
<GID>36</GID>
<name>ENABLE_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-29,76.5,-29</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-37,68,-32.5</points>
<connection>
<GID>41</GID>
<name>OUT_2</name></connection>
<connection>
<GID>36</GID>
<name>DATA_IN_2</name></connection>
<connection>
<GID>36</GID>
<name>DATA_OUT_2</name></connection>
<intersection>-34.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>56,-34.5,68,-34.5</points>
<intersection>56 9</intersection>
<intersection>68 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>56,-43,56,-34.5</points>
<connection>
<GID>47</GID>
<name>N_in3</name></connection>
<intersection>-34.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-37,69,-32.5</points>
<connection>
<GID>41</GID>
<name>OUT_1</name></connection>
<connection>
<GID>36</GID>
<name>DATA_IN_1</name></connection>
<connection>
<GID>36</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-35 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>58.5,-35,69,-35</points>
<intersection>58.5 9</intersection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>58.5,-43,58.5,-35</points>
<connection>
<GID>48</GID>
<name>N_in3</name></connection>
<intersection>-35 8</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-37,70,-32.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<connection>
<GID>36</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>36</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-35.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>61,-35.5,70,-35.5</points>
<intersection>61 9</intersection>
<intersection>70 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>61,-43,61,-35.5</points>
<connection>
<GID>49</GID>
<name>N_in3</name></connection>
<intersection>-35.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-37,67,-32.5</points>
<connection>
<GID>41</GID>
<name>OUT_3</name></connection>
<connection>
<GID>36</GID>
<name>DATA_IN_3</name></connection>
<connection>
<GID>36</GID>
<name>DATA_OUT_3</name></connection>
<intersection>-34 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>53.5,-34,67,-34</points>
<intersection>53.5 9</intersection>
<intersection>67 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>53.5,-43,53.5,-34</points>
<connection>
<GID>46</GID>
<name>N_in3</name></connection>
<intersection>-34 8</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-46.5,71.5,-43.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-43.5,70,-41</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-43.5,71.5,-43.5</points>
<intersection>70 1</intersection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-46.5,69.5,-43.5</points>
<connection>
<GID>51</GID>
<name>OUT_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>69,-43.5,69,-41</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-43.5,69.5,-43.5</points>
<intersection>69 1</intersection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-46.5,67.5,-43.5</points>
<connection>
<GID>51</GID>
<name>OUT_2</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68,-43.5,68,-41</points>
<connection>
<GID>41</GID>
<name>IN_2</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-43.5,68,-43.5</points>
<intersection>67.5 0</intersection>
<intersection>68 1</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-46.5,65.5,-43.5</points>
<connection>
<GID>51</GID>
<name>OUT_3</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>67,-43.5,67,-41</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-43.5,67,-43.5</points>
<intersection>65.5 0</intersection>
<intersection>67 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-50,53.5,-45</points>
<connection>
<GID>46</GID>
<name>N_in2</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-50,55.5,-50</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-53,55,-46.5</points>
<intersection>-53 4</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-46.5,61,-46.5</points>
<intersection>55 0</intersection>
<intersection>61 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>61,-46.5,61,-45</points>
<connection>
<GID>49</GID>
<name>N_in2</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>55,-53,55.5,-53</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-51,54,-45.5</points>
<intersection>-51 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-51,55.5,-51</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-45.5,56,-45.5</points>
<intersection>54 0</intersection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-45.5,56,-45</points>
<connection>
<GID>47</GID>
<name>N_in2</name></connection>
<intersection>-45.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-52,54.5,-46</points>
<intersection>-52 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-52,55.5,-52</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-46,58.5,-46</points>
<intersection>54.5 0</intersection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-46,58.5,-45</points>
<connection>
<GID>48</GID>
<name>N_in2</name></connection>
<intersection>-46 2</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>