<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>493.5,1544.74,775.175,1360.77</PageViewport>
<gate>
<ID>1538</ID>
<type>DE_TO</type>
<position>758.5,1435.5</position>
<input>
<ID>IN_0</ID>1719 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>1539</ID>
<type>DE_TO</type>
<position>763.5,1436.5</position>
<input>
<ID>IN_0</ID>1718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>1540</ID>
<type>DE_TO</type>
<position>758.5,1437.5</position>
<input>
<ID>IN_0</ID>1717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>2</ID>
<type>AM_REGISTER16</type>
<position>512.5,1507.5</position>
<input>
<ID>clear</ID>4 </input>
<input>
<ID>clock</ID>5 </input>
<input>
<ID>count_enable</ID>8 </input>
<input>
<ID>count_up</ID>3 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1541</ID>
<type>DE_TO</type>
<position>763.5,1438.5</position>
<input>
<ID>IN_0</ID>1716 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>3</ID>
<type>BA_NAND4</type>
<position>728,1504</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>1611 </input>
<input>
<ID>IN_2</ID>1610 </input>
<input>
<ID>IN_3</ID>1609 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1542</ID>
<type>BA_NAND3</type>
<position>751.5,1447.5</position>
<input>
<ID>IN_0</ID>1721 </input>
<input>
<ID>IN_1</ID>1722 </input>
<input>
<ID>IN_2</ID>1723 </input>
<output>
<ID>OUT</ID>1720 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>513.5,1523</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1543</ID>
<type>DA_FROM</type>
<position>753.5,1454.5</position>
<input>
<ID>IN_0</ID>1721 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID OC0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>519.5,1520.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1544</ID>
<type>DA_FROM</type>
<position>751.5,1454.5</position>
<input>
<ID>IN_0</ID>1722 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID OC1</lparam></gate>
<gate>
<ID>6</ID>
<type>EE_VDD</type>
<position>524,1522.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1545</ID>
<type>AE_OR2</type>
<position>595,1390</position>
<input>
<ID>IN_0</ID>1619 </input>
<input>
<ID>IN_1</ID>1617 </input>
<output>
<ID>OUT</ID>1614 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>734.5,1499</position>
<input>
<ID>IN_0</ID>1612 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1546</ID>
<type>DA_FROM</type>
<position>749.5,1454.5</position>
<input>
<ID>IN_0</ID>1723 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID OC2</lparam></gate>
<gate>
<ID>1547</ID>
<type>AE_OR2</type>
<position>550.5,1411.5</position>
<input>
<ID>IN_0</ID>1738 </input>
<input>
<ID>IN_1</ID>1739 </input>
<output>
<ID>OUT</ID>1737 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>506,1485.5</position>
<gparam>LABEL_TEXT RESET LICZNIKA</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1548</ID>
<type>AA_AND2</type>
<position>744,1431.5</position>
<input>
<ID>IN_0</ID>1720 </input>
<input>
<ID>IN_1</ID>1743 </input>
<output>
<ID>OUT</ID>1724 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>529,1505.5</position>
<input>
<ID>IN_0</ID>1392 </input>
<input>
<ID>IN_1</ID>1389 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1549</ID>
<type>CC_PULSE</type>
<position>543.5,1412.5</position>
<output>
<ID>OUT_0</ID>1738 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1550</ID>
<type>DA_FROM</type>
<position>579.5,1394</position>
<input>
<ID>IN_0</ID>1620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW3</lparam></gate>
<gate>
<ID>12</ID>
<type>CC_PULSE</type>
<position>506,1488</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1551</ID>
<type>DA_FROM</type>
<position>755,1422</position>
<input>
<ID>IN_0</ID>1745 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>515.5,1526</position>
<gparam>LABEL_TEXT LICZNIK ON OFF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1552</ID>
<type>DA_FROM</type>
<position>538,1410.5</position>
<input>
<ID>IN_0</ID>1739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Do step</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR2</type>
<position>511.5,1494</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1553</ID>
<type>DA_FROM</type>
<position>752.5,1424</position>
<input>
<ID>IN_0</ID>1744 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1554</ID>
<type>DA_FROM</type>
<position>585.5,1384</position>
<input>
<ID>IN_0</ID>1617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1555</ID>
<type>AA_LABEL</type>
<position>544.5,1415.5</position>
<gparam>LABEL_TEXT step</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1556</ID>
<type>AE_OR2</type>
<position>761,1429</position>
<input>
<ID>IN_0</ID>1727 </input>
<input>
<ID>IN_1</ID>1726 </input>
<output>
<ID>OUT</ID>1725 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1557</ID>
<type>AE_OR4</type>
<position>584.5,1391</position>
<input>
<ID>IN_0</ID>1620 </input>
<input>
<ID>IN_1</ID>1621 </input>
<input>
<ID>IN_2</ID>1622 </input>
<input>
<ID>IN_3</ID>1623 </input>
<output>
<ID>OUT</ID>1619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1558</ID>
<type>DA_FROM</type>
<position>579.5,1392</position>
<input>
<ID>IN_0</ID>1621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW2</lparam></gate>
<gate>
<ID>1559</ID>
<type>DA_FROM</type>
<position>579.5,1390</position>
<input>
<ID>IN_0</ID>1622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW1</lparam></gate>
<gate>
<ID>1560</ID>
<type>DA_FROM</type>
<position>578,1388</position>
<input>
<ID>IN_0</ID>1623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW</lparam></gate>
<gate>
<ID>1561</ID>
<type>DA_FROM</type>
<position>770.5,1430.5</position>
<input>
<ID>IN_0</ID>1726 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID TCR</lparam></gate>
<gate>
<ID>1562</ID>
<type>AM_RAM_16x16</type>
<position>669,1428.5</position>
<input>
<ID>ADDRESS_0</ID>1624 </input>
<input>
<ID>ADDRESS_1</ID>1625 </input>
<input>
<ID>ADDRESS_10</ID>1634 </input>
<input>
<ID>ADDRESS_11</ID>1635 </input>
<input>
<ID>ADDRESS_12</ID>1636 </input>
<input>
<ID>ADDRESS_13</ID>1637 </input>
<input>
<ID>ADDRESS_14</ID>1638 </input>
<input>
<ID>ADDRESS_15</ID>1639 </input>
<input>
<ID>ADDRESS_2</ID>1626 </input>
<input>
<ID>ADDRESS_3</ID>1627 </input>
<input>
<ID>ADDRESS_4</ID>1628 </input>
<input>
<ID>ADDRESS_5</ID>1629 </input>
<input>
<ID>ADDRESS_6</ID>1630 </input>
<input>
<ID>ADDRESS_7</ID>1631 </input>
<input>
<ID>ADDRESS_8</ID>1632 </input>
<input>
<ID>ADDRESS_9</ID>1633 </input>
<input>
<ID>DATA_IN_0</ID>1643 </input>
<input>
<ID>DATA_IN_1</ID>1644 </input>
<input>
<ID>DATA_IN_10</ID>1653 </input>
<input>
<ID>DATA_IN_11</ID>1654 </input>
<input>
<ID>DATA_IN_12</ID>1655 </input>
<input>
<ID>DATA_IN_13</ID>1656 </input>
<input>
<ID>DATA_IN_14</ID>1657 </input>
<input>
<ID>DATA_IN_15</ID>1658 </input>
<input>
<ID>DATA_IN_2</ID>1645 </input>
<input>
<ID>DATA_IN_3</ID>1646 </input>
<input>
<ID>DATA_IN_4</ID>1647 </input>
<input>
<ID>DATA_IN_5</ID>1648 </input>
<input>
<ID>DATA_IN_6</ID>1649 </input>
<input>
<ID>DATA_IN_7</ID>1650 </input>
<input>
<ID>DATA_IN_8</ID>1651 </input>
<input>
<ID>DATA_IN_9</ID>1652 </input>
<output>
<ID>DATA_OUT_0</ID>1643 </output>
<output>
<ID>DATA_OUT_1</ID>1644 </output>
<output>
<ID>DATA_OUT_10</ID>1653 </output>
<output>
<ID>DATA_OUT_11</ID>1654 </output>
<output>
<ID>DATA_OUT_12</ID>1655 </output>
<output>
<ID>DATA_OUT_13</ID>1656 </output>
<output>
<ID>DATA_OUT_14</ID>1657 </output>
<output>
<ID>DATA_OUT_15</ID>1658 </output>
<output>
<ID>DATA_OUT_2</ID>1645 </output>
<output>
<ID>DATA_OUT_3</ID>1646 </output>
<output>
<ID>DATA_OUT_4</ID>1647 </output>
<output>
<ID>DATA_OUT_5</ID>1648 </output>
<output>
<ID>DATA_OUT_6</ID>1649 </output>
<output>
<ID>DATA_OUT_7</ID>1650 </output>
<output>
<ID>DATA_OUT_8</ID>1651 </output>
<output>
<ID>DATA_OUT_9</ID>1652 </output>
<input>
<ID>ENABLE_0</ID>1359 </input>
<input>
<ID>write_clock</ID>1616 </input>
<input>
<ID>write_enable</ID>1360 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 16</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 6144</lparam>
<lparam>Address:1 14338</lparam>
<lparam>Address:2 10241</lparam>
<lparam>Address:3 28672</lparam>
<lparam>Address:2048 65534</lparam>
<lparam>Address:2050 1</lparam></gate>
<gate>
<ID>1563</ID>
<type>DA_FROM</type>
<position>767,1427.5</position>
<input>
<ID>IN_0</ID>1727 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1564</ID>
<type>AM_REGISTER16</type>
<position>650.5,1428.5</position>
<input>
<ID>IN_0</ID>1409 </input>
<input>
<ID>IN_1</ID>1400 </input>
<input>
<ID>IN_10</ID>1412 </input>
<input>
<ID>IN_11</ID>1404 </input>
<input>
<ID>IN_12</ID>1411 </input>
<input>
<ID>IN_13</ID>1403 </input>
<input>
<ID>IN_14</ID>1410 </input>
<input>
<ID>IN_15</ID>1402 </input>
<input>
<ID>IN_2</ID>1408 </input>
<input>
<ID>IN_3</ID>1401 </input>
<input>
<ID>IN_4</ID>1415 </input>
<input>
<ID>IN_5</ID>1407 </input>
<input>
<ID>IN_6</ID>1414 </input>
<input>
<ID>IN_7</ID>1406 </input>
<input>
<ID>IN_8</ID>1413 </input>
<input>
<ID>IN_9</ID>1405 </input>
<output>
<ID>OUT_0</ID>1624 </output>
<output>
<ID>OUT_1</ID>1625 </output>
<output>
<ID>OUT_10</ID>1634 </output>
<output>
<ID>OUT_11</ID>1635 </output>
<output>
<ID>OUT_12</ID>1636 </output>
<output>
<ID>OUT_13</ID>1637 </output>
<output>
<ID>OUT_14</ID>1638 </output>
<output>
<ID>OUT_15</ID>1639 </output>
<output>
<ID>OUT_2</ID>1626 </output>
<output>
<ID>OUT_3</ID>1627 </output>
<output>
<ID>OUT_4</ID>1628 </output>
<output>
<ID>OUT_5</ID>1629 </output>
<output>
<ID>OUT_6</ID>1630 </output>
<output>
<ID>OUT_7</ID>1631 </output>
<output>
<ID>OUT_8</ID>1632 </output>
<output>
<ID>OUT_9</ID>1633 </output>
<input>
<ID>clear</ID>1691 </input>
<input>
<ID>clock</ID>1640 </input>
<input>
<ID>load</ID>1491 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1565</ID>
<type>AA_AND2</type>
<position>553.5,1430</position>
<input>
<ID>IN_0</ID>1736 </input>
<input>
<ID>IN_1</ID>1730 </input>
<output>
<ID>OUT</ID>1728 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1566</ID>
<type>AE_OR2</type>
<position>646,1416.5</position>
<input>
<ID>IN_0</ID>1641 </input>
<input>
<ID>IN_1</ID>1642 </input>
<output>
<ID>OUT</ID>1640 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1567</ID>
<type>AE_OR2</type>
<position>564,1429</position>
<input>
<ID>IN_0</ID>1728 </input>
<input>
<ID>IN_1</ID>1729 </input>
<output>
<ID>OUT</ID>1731 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1568</ID>
<type>DA_FROM</type>
<position>638,1417.5</position>
<input>
<ID>IN_0</ID>1641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MARW</lparam></gate>
<gate>
<ID>1569</ID>
<type>DA_FROM</type>
<position>641,1415.5</position>
<input>
<ID>IN_0</ID>1642 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1570</ID>
<type>AE_SMALL_INVERTER</type>
<position>557,1426.5</position>
<input>
<ID>IN_0</ID>1730 </input>
<output>
<ID>OUT_0</ID>1729 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1571</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>668.5,1406.5</position>
<input>
<ID>ENABLE_0</ID>1359 </input>
<input>
<ID>IN_0</ID>1658 </input>
<input>
<ID>IN_1</ID>1657 </input>
<input>
<ID>IN_10</ID>1648 </input>
<input>
<ID>IN_11</ID>1647 </input>
<input>
<ID>IN_12</ID>1646 </input>
<input>
<ID>IN_13</ID>1645 </input>
<input>
<ID>IN_14</ID>1644 </input>
<input>
<ID>IN_15</ID>1643 </input>
<input>
<ID>IN_2</ID>1656 </input>
<input>
<ID>IN_3</ID>1655 </input>
<input>
<ID>IN_4</ID>1654 </input>
<input>
<ID>IN_5</ID>1653 </input>
<input>
<ID>IN_6</ID>1652 </input>
<input>
<ID>IN_7</ID>1651 </input>
<input>
<ID>IN_8</ID>1650 </input>
<input>
<ID>IN_9</ID>1649 </input>
<output>
<ID>OUT_0</ID>1666 </output>
<output>
<ID>OUT_1</ID>1683 </output>
<output>
<ID>OUT_10</ID>1661 </output>
<output>
<ID>OUT_11</ID>1688 </output>
<output>
<ID>OUT_12</ID>1660 </output>
<output>
<ID>OUT_13</ID>1689 </output>
<output>
<ID>OUT_14</ID>1659 </output>
<output>
<ID>OUT_15</ID>1690 </output>
<output>
<ID>OUT_2</ID>1665 </output>
<output>
<ID>OUT_3</ID>1684 </output>
<output>
<ID>OUT_4</ID>1664 </output>
<output>
<ID>OUT_5</ID>1685 </output>
<output>
<ID>OUT_6</ID>1663 </output>
<output>
<ID>OUT_7</ID>1686 </output>
<output>
<ID>OUT_8</ID>1662 </output>
<output>
<ID>OUT_9</ID>1687 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1572</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>695.5,1406</position>
<input>
<ID>ENABLE_0</ID>1360 </input>
<input>
<ID>IN_0</ID>1675 </input>
<input>
<ID>IN_1</ID>1674 </input>
<input>
<ID>IN_10</ID>1680 </input>
<input>
<ID>IN_11</ID>1668 </input>
<input>
<ID>IN_12</ID>1681 </input>
<input>
<ID>IN_13</ID>1669 </input>
<input>
<ID>IN_14</ID>1682 </input>
<input>
<ID>IN_15</ID>1667 </input>
<input>
<ID>IN_2</ID>1676 </input>
<input>
<ID>IN_3</ID>1673 </input>
<input>
<ID>IN_4</ID>1677 </input>
<input>
<ID>IN_5</ID>1672 </input>
<input>
<ID>IN_6</ID>1678 </input>
<input>
<ID>IN_7</ID>1671 </input>
<input>
<ID>IN_8</ID>1679 </input>
<input>
<ID>IN_9</ID>1670 </input>
<output>
<ID>OUT_0</ID>1643 </output>
<output>
<ID>OUT_1</ID>1644 </output>
<output>
<ID>OUT_10</ID>1653 </output>
<output>
<ID>OUT_11</ID>1654 </output>
<output>
<ID>OUT_12</ID>1655 </output>
<output>
<ID>OUT_13</ID>1656 </output>
<output>
<ID>OUT_14</ID>1657 </output>
<output>
<ID>OUT_15</ID>1658 </output>
<output>
<ID>OUT_2</ID>1645 </output>
<output>
<ID>OUT_3</ID>1646 </output>
<output>
<ID>OUT_4</ID>1647 </output>
<output>
<ID>OUT_5</ID>1648 </output>
<output>
<ID>OUT_6</ID>1649 </output>
<output>
<ID>OUT_7</ID>1650 </output>
<output>
<ID>OUT_8</ID>1651 </output>
<output>
<ID>OUT_9</ID>1652 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1573</ID>
<type>DE_TO</type>
<position>661,1394.5</position>
<input>
<ID>IN_0</ID>1666 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1574</ID>
<type>DE_TO</type>
<position>663,1394.5</position>
<input>
<ID>IN_0</ID>1665 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1575</ID>
<type>DE_TO</type>
<position>665,1394.5</position>
<input>
<ID>IN_0</ID>1664 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1576</ID>
<type>DE_TO</type>
<position>667,1394.5</position>
<input>
<ID>IN_0</ID>1663 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1577</ID>
<type>DE_TO</type>
<position>669,1394.5</position>
<input>
<ID>IN_0</ID>1662 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1578</ID>
<type>DE_TO</type>
<position>671,1394.5</position>
<input>
<ID>IN_0</ID>1661 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1579</ID>
<type>DE_TO</type>
<position>673,1394.5</position>
<input>
<ID>IN_0</ID>1660 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1580</ID>
<type>DE_TO</type>
<position>675,1394.5</position>
<input>
<ID>IN_0</ID>1659 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1581</ID>
<type>DE_TO</type>
<position>688,1392</position>
<input>
<ID>IN_0</ID>1667 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1582</ID>
<type>DE_TO</type>
<position>690,1392</position>
<input>
<ID>IN_0</ID>1669 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1583</ID>
<type>DE_TO</type>
<position>692,1392</position>
<input>
<ID>IN_0</ID>1668 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1584</ID>
<type>DE_TO</type>
<position>694,1392</position>
<input>
<ID>IN_0</ID>1670 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1585</ID>
<type>DE_TO</type>
<position>696,1392</position>
<input>
<ID>IN_0</ID>1671 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1586</ID>
<type>DE_TO</type>
<position>698,1392</position>
<input>
<ID>IN_0</ID>1672 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1587</ID>
<type>DE_TO</type>
<position>700,1392</position>
<input>
<ID>IN_0</ID>1673 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1588</ID>
<type>DE_TO</type>
<position>702,1392</position>
<input>
<ID>IN_0</ID>1674 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1589</ID>
<type>DE_TO</type>
<position>689,1399.5</position>
<input>
<ID>IN_0</ID>1682 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1590</ID>
<type>DE_TO</type>
<position>691,1399.5</position>
<input>
<ID>IN_0</ID>1681 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1591</ID>
<type>DE_TO</type>
<position>693,1399.5</position>
<input>
<ID>IN_0</ID>1680 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1592</ID>
<type>DE_TO</type>
<position>695,1399.5</position>
<input>
<ID>IN_0</ID>1679 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1593</ID>
<type>DE_TO</type>
<position>697,1399.5</position>
<input>
<ID>IN_0</ID>1678 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1594</ID>
<type>DE_TO</type>
<position>699,1399.5</position>
<input>
<ID>IN_0</ID>1677 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1595</ID>
<type>DE_TO</type>
<position>701,1399.5</position>
<input>
<ID>IN_0</ID>1676 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1596</ID>
<type>DE_TO</type>
<position>703,1399.5</position>
<input>
<ID>IN_0</ID>1675 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1597</ID>
<type>DE_TO</type>
<position>662,1401.5</position>
<input>
<ID>IN_0</ID>1683 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1598</ID>
<type>DE_TO</type>
<position>664,1401.5</position>
<input>
<ID>IN_0</ID>1684 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1599</ID>
<type>DE_TO</type>
<position>666,1401.5</position>
<input>
<ID>IN_0</ID>1685 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1600</ID>
<type>DE_TO</type>
<position>668,1401.5</position>
<input>
<ID>IN_0</ID>1686 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1601</ID>
<type>DE_TO</type>
<position>670,1401.5</position>
<input>
<ID>IN_0</ID>1687 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1602</ID>
<type>DE_TO</type>
<position>672,1401.5</position>
<input>
<ID>IN_0</ID>1688 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1603</ID>
<type>DE_TO</type>
<position>674,1401.5</position>
<input>
<ID>IN_0</ID>1689 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1604</ID>
<type>DE_TO</type>
<position>676,1401.5</position>
<input>
<ID>IN_0</ID>1690 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1605</ID>
<type>DE_TO</type>
<position>577.5,1422</position>
<input>
<ID>IN_0</ID>1732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>1606</ID>
<type>DA_FROM</type>
<position>654.5,1415.5</position>
<input>
<ID>IN_0</ID>1691 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1607</ID>
<type>AA_AND2</type>
<position>570.5,1422</position>
<input>
<ID>IN_0</ID>1731 </input>
<input>
<ID>IN_1</ID>1733 </input>
<output>
<ID>OUT</ID>1732 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1608</ID>
<type>DA_FROM</type>
<position>685,1402</position>
<input>
<ID>IN_0</ID>1360 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ACS</lparam></gate>
<gate>
<ID>1609</ID>
<type>AE_OR2</type>
<position>562.5,1421</position>
<input>
<ID>IN_0</ID>1734 </input>
<input>
<ID>IN_1</ID>1737 </input>
<output>
<ID>OUT</ID>1733 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1610</ID>
<type>AA_AND2</type>
<position>553.5,1422</position>
<input>
<ID>IN_0</ID>1361 </input>
<input>
<ID>IN_1</ID>1735 </input>
<output>
<ID>OUT</ID>1734 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1611</ID>
<type>AE_OR2</type>
<position>745.5,1423</position>
<input>
<ID>IN_0</ID>1745 </input>
<input>
<ID>IN_1</ID>1744 </input>
<output>
<ID>OUT</ID>1743 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1612</ID>
<type>FF_GND</type>
<position>717.5,1445.5</position>
<output>
<ID>OUT_0</ID>1740 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1613</ID>
<type>DA_FROM</type>
<position>545,1421</position>
<input>
<ID>IN_0</ID>1735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Start</lparam></gate>
<gate>
<ID>1614</ID>
<type>EE_VDD</type>
<position>738,1439</position>
<output>
<ID>OUT_0</ID>1741 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1615</ID>
<type>DA_FROM</type>
<position>542.5,1431</position>
<input>
<ID>IN_0</ID>1736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input</lparam></gate>
<gate>
<ID>1616</ID>
<type>DA_FROM</type>
<position>545,1428</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InS</lparam></gate>
<gate>
<ID>1617</ID>
<type>DE_TO</type>
<position>737,1419</position>
<input>
<ID>IN_0</ID>1692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TCR</lparam></gate>
<gate>
<ID>1618</ID>
<type>DE_TO</type>
<position>737,1417</position>
<input>
<ID>IN_0</ID>1693 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALUS</lparam></gate>
<gate>
<ID>1619</ID>
<type>AA_LABEL</type>
<position>723,1450</position>
<gparam>LABEL_TEXT Control Unite</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1620</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>575.5,1470.5</position>
<input>
<ID>ENABLE_0</ID>1341 </input>
<input>
<ID>IN_0</ID>1380 </input>
<input>
<ID>IN_1</ID>1387 </input>
<input>
<ID>IN_10</ID>1384 </input>
<input>
<ID>IN_12</ID>1385 </input>
<input>
<ID>IN_14</ID>1386 </input>
<input>
<ID>IN_15</ID>1388 </input>
<input>
<ID>IN_2</ID>1381 </input>
<input>
<ID>IN_4</ID>1379 </input>
<input>
<ID>IN_6</ID>1382 </input>
<input>
<ID>IN_8</ID>1383 </input>
<output>
<ID>OUT_0</ID>1762 </output>
<output>
<ID>OUT_1</ID>1763 </output>
<output>
<ID>OUT_10</ID>1772 </output>
<output>
<ID>OUT_11</ID>1773 </output>
<output>
<ID>OUT_12</ID>1774 </output>
<output>
<ID>OUT_13</ID>1775 </output>
<output>
<ID>OUT_14</ID>1776 </output>
<output>
<ID>OUT_15</ID>1777 </output>
<output>
<ID>OUT_2</ID>1764 </output>
<output>
<ID>OUT_3</ID>1765 </output>
<output>
<ID>OUT_4</ID>1766 </output>
<output>
<ID>OUT_5</ID>1767 </output>
<output>
<ID>OUT_6</ID>1768 </output>
<output>
<ID>OUT_7</ID>1769 </output>
<output>
<ID>OUT_8</ID>1770 </output>
<output>
<ID>OUT_9</ID>1771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1621</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>564.5,1449.5</position>
<input>
<ID>ENABLE_0</ID>1778 </input>
<input>
<ID>IN_0</ID>1757 </input>
<input>
<ID>IN_1</ID>1753 </input>
<input>
<ID>IN_10</ID>1760 </input>
<input>
<ID>IN_11</ID>1748 </input>
<input>
<ID>IN_12</ID>1759 </input>
<input>
<ID>IN_13</ID>1747 </input>
<input>
<ID>IN_14</ID>1758 </input>
<input>
<ID>IN_15</ID>1746 </input>
<input>
<ID>IN_2</ID>1756 </input>
<input>
<ID>IN_3</ID>1752 </input>
<input>
<ID>IN_4</ID>1755 </input>
<input>
<ID>IN_5</ID>1751 </input>
<input>
<ID>IN_6</ID>1754 </input>
<input>
<ID>IN_7</ID>1750 </input>
<input>
<ID>IN_8</ID>1761 </input>
<input>
<ID>IN_9</ID>1749 </input>
<output>
<ID>OUT_0</ID>1762 </output>
<output>
<ID>OUT_1</ID>1763 </output>
<output>
<ID>OUT_10</ID>1772 </output>
<output>
<ID>OUT_11</ID>1773 </output>
<output>
<ID>OUT_12</ID>1774 </output>
<output>
<ID>OUT_13</ID>1775 </output>
<output>
<ID>OUT_14</ID>1776 </output>
<output>
<ID>OUT_15</ID>1777 </output>
<output>
<ID>OUT_2</ID>1764 </output>
<output>
<ID>OUT_3</ID>1765 </output>
<output>
<ID>OUT_4</ID>1766 </output>
<output>
<ID>OUT_5</ID>1767 </output>
<output>
<ID>OUT_6</ID>1768 </output>
<output>
<ID>OUT_7</ID>1769 </output>
<output>
<ID>OUT_8</ID>1770 </output>
<output>
<ID>OUT_9</ID>1771 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1622</ID>
<type>AA_TOGGLE</type>
<position>559,1460.5</position>
<output>
<ID>OUT_0</ID>1778 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1195</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>621,1475.5</position>
<input>
<ID>ENABLE_0</ID>1373 </input>
<input>
<ID>IN_0</ID>1432 </input>
<input>
<ID>IN_1</ID>1424 </input>
<input>
<ID>IN_10</ID>1427 </input>
<input>
<ID>IN_11</ID>1420 </input>
<input>
<ID>IN_12</ID>1426 </input>
<input>
<ID>IN_13</ID>1419 </input>
<input>
<ID>IN_14</ID>1425 </input>
<input>
<ID>IN_15</ID>1418 </input>
<input>
<ID>IN_2</ID>1431 </input>
<input>
<ID>IN_3</ID>1423 </input>
<input>
<ID>IN_4</ID>1430 </input>
<input>
<ID>IN_5</ID>1422 </input>
<input>
<ID>IN_6</ID>1429 </input>
<input>
<ID>IN_7</ID>1421 </input>
<input>
<ID>IN_8</ID>1428 </input>
<input>
<ID>IN_9</ID>1417 </input>
<output>
<ID>OUT_0</ID>1336 </output>
<output>
<ID>OUT_1</ID>1328 </output>
<output>
<ID>OUT_10</ID>1331 </output>
<output>
<ID>OUT_11</ID>1323 </output>
<output>
<ID>OUT_12</ID>1330 </output>
<output>
<ID>OUT_13</ID>1322 </output>
<output>
<ID>OUT_14</ID>1329 </output>
<output>
<ID>OUT_15</ID>1321 </output>
<output>
<ID>OUT_2</ID>1335 </output>
<output>
<ID>OUT_3</ID>1327 </output>
<output>
<ID>OUT_4</ID>1334 </output>
<output>
<ID>OUT_5</ID>1326 </output>
<output>
<ID>OUT_6</ID>1333 </output>
<output>
<ID>OUT_7</ID>1325 </output>
<output>
<ID>OUT_8</ID>1332 </output>
<output>
<ID>OUT_9</ID>1324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1196</ID>
<type>GA_LED</type>
<position>537,1490.5</position>
<input>
<ID>N_in0</ID>1337 </input>
<input>
<ID>N_in1</ID>1338 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1197</ID>
<type>BI_DECODER_4x16</type>
<position>522,1473.5</position>
<input>
<ID>ENABLE</ID>1353 </input>
<input>
<ID>IN_0</ID>1357 </input>
<input>
<ID>IN_1</ID>1356 </input>
<input>
<ID>IN_2</ID>1355 </input>
<input>
<ID>IN_3</ID>1354 </input>
<output>
<ID>OUT_0</ID>1339 </output>
<output>
<ID>OUT_1</ID>1340 </output>
<output>
<ID>OUT_11</ID>1372 </output>
<output>
<ID>OUT_13</ID>1391 </output>
<output>
<ID>OUT_2</ID>1347 </output>
<output>
<ID>OUT_3</ID>1349 </output>
<output>
<ID>OUT_4</ID>1363 </output>
<output>
<ID>OUT_5</ID>1351 </output>
<output>
<ID>OUT_6</ID>1352 </output>
<output>
<ID>OUT_8</ID>1337 </output>
<output>
<ID>OUT_9</ID>1358 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1198</ID>
<type>DA_FROM</type>
<position>651.5,1487</position>
<input>
<ID>IN_0</ID>1376 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Add X</lparam></gate>
<gate>
<ID>1199</ID>
<type>AA_TOGGLE</type>
<position>528,1434.5</position>
<output>
<ID>OUT_0</ID>1730 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1200</ID>
<type>DE_TO</type>
<position>542,1466</position>
<input>
<ID>IN_0</ID>1340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Load X</lparam></gate>
<gate>
<ID>1201</ID>
<type>DE_TO</type>
<position>542,1469</position>
<input>
<ID>IN_0</ID>1347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Store X</lparam></gate>
<gate>
<ID>1202</ID>
<type>AE_OR4</type>
<position>643,1488</position>
<input>
<ID>IN_0</ID>1377 </input>
<input>
<ID>IN_1</ID>1376 </input>
<input>
<ID>IN_2</ID>1375 </input>
<input>
<ID>IN_3</ID>1396 </input>
<output>
<ID>OUT</ID>1373 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1203</ID>
<type>DA_FROM</type>
<position>659.5,1496.5</position>
<input>
<ID>IN_0</ID>1394 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AddI X</lparam></gate>
<gate>
<ID>1204</ID>
<type>CC_PULSE</type>
<position>533,1425</position>
<output>
<ID>OUT_0</ID>1361 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1205</ID>
<type>DA_FROM</type>
<position>651.5,1484.5</position>
<input>
<ID>IN_0</ID>1377 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Subt X</lparam></gate>
<gate>
<ID>1206</ID>
<type>BB_CLOCK</type>
<position>553,1500.5</position>
<output>
<ID>CLK</ID>1397 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>1207</ID>
<type>AA_LABEL</type>
<position>541.5,1519.5</position>
<gparam>LABEL_TEXT 1-start/0-stop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1208</ID>
<type>AA_AND2</type>
<position>581.5,1506.5</position>
<input>
<ID>IN_0</ID>1389 </input>
<input>
<ID>IN_1</ID>1392 </input>
<output>
<ID>OUT</ID>1573 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1209</ID>
<type>AA_TOGGLE</type>
<position>555.5,1518.5</position>
<output>
<ID>OUT_0</ID>1389 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1210</ID>
<type>DA_FROM</type>
<position>701.5,1496</position>
<input>
<ID>IN_0</ID>1342 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1211</ID>
<type>DE_TO</type>
<position>747,1496.5</position>
<input>
<ID>IN_0</ID>1576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>1212</ID>
<type>DE_TO</type>
<position>747,1494</position>
<input>
<ID>IN_0</ID>1581 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>1213</ID>
<type>DA_FROM</type>
<position>701.5,1494</position>
<input>
<ID>IN_0</ID>1343 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1214</ID>
<type>AA_LABEL</type>
<position>763.5,1487</position>
<gparam>LABEL_TEXT KOD ROZKAZU</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1215</ID>
<type>DA_FROM</type>
<position>701.5,1492</position>
<input>
<ID>IN_0</ID>1344 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1216</ID>
<type>AA_LABEL</type>
<position>752,1499.5</position>
<gparam>LABEL_TEXT WARUNKI SKOKU</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1217</ID>
<type>DA_FROM</type>
<position>701.5,1490</position>
<input>
<ID>IN_0</ID>1345 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1218</ID>
<type>DE_TO</type>
<position>542,1472</position>
<input>
<ID>IN_0</ID>1349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Add X</lparam></gate>
<gate>
<ID>1219</ID>
<type>CC_PULSE</type>
<position>556.5,1510.5</position>
<output>
<ID>OUT_0</ID>1390 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1220</ID>
<type>AE_OR2</type>
<position>650,1496</position>
<input>
<ID>IN_0</ID>1395 </input>
<input>
<ID>IN_1</ID>1394 </input>
<output>
<ID>OUT</ID>1396 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1221</ID>
<type>DE_TO</type>
<position>657,1493</position>
<input>
<ID>IN_0</ID>1395 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond1</lparam></gate>
<gate>
<ID>1222</ID>
<type>DE_TO</type>
<position>543,1499</position>
<input>
<ID>IN_0</ID>1391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LoadI</lparam></gate>
<gate>
<ID>1223</ID>
<type>DE_TO</type>
<position>635,1506</position>
<input>
<ID>IN_0</ID>1418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k15</lparam></gate>
<gate>
<ID>1224</ID>
<type>DE_TO</type>
<position>635,1504</position>
<input>
<ID>IN_0</ID>1419 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k13</lparam></gate>
<gate>
<ID>1225</ID>
<type>DE_TO</type>
<position>635,1502</position>
<input>
<ID>IN_0</ID>1420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k11</lparam></gate>
<gate>
<ID>1226</ID>
<type>DE_TO</type>
<position>635,1500</position>
<input>
<ID>IN_0</ID>1417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k9</lparam></gate>
<gate>
<ID>1227</ID>
<type>DE_TO</type>
<position>635,1498</position>
<input>
<ID>IN_0</ID>1421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k7</lparam></gate>
<gate>
<ID>1228</ID>
<type>DE_TO</type>
<position>635,1496</position>
<input>
<ID>IN_0</ID>1422 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k5</lparam></gate>
<gate>
<ID>1229</ID>
<type>DE_TO</type>
<position>635,1494</position>
<input>
<ID>IN_0</ID>1423 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k3</lparam></gate>
<gate>
<ID>1230</ID>
<type>DE_TO</type>
<position>635,1492</position>
<input>
<ID>IN_0</ID>1424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k1</lparam></gate>
<gate>
<ID>1231</ID>
<type>DE_TO</type>
<position>628,1505</position>
<input>
<ID>IN_0</ID>1425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k14</lparam></gate>
<gate>
<ID>1232</ID>
<type>DE_TO</type>
<position>628,1503</position>
<input>
<ID>IN_0</ID>1426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k12</lparam></gate>
<gate>
<ID>1233</ID>
<type>DE_TO</type>
<position>628,1501</position>
<input>
<ID>IN_0</ID>1427 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k10</lparam></gate>
<gate>
<ID>1234</ID>
<type>DE_TO</type>
<position>628,1499</position>
<input>
<ID>IN_0</ID>1428 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k8</lparam></gate>
<gate>
<ID>1235</ID>
<type>DE_TO</type>
<position>628,1497</position>
<input>
<ID>IN_0</ID>1429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k6</lparam></gate>
<gate>
<ID>1236</ID>
<type>DE_TO</type>
<position>628,1495</position>
<input>
<ID>IN_0</ID>1430 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k4</lparam></gate>
<gate>
<ID>1237</ID>
<type>DE_TO</type>
<position>628,1493</position>
<input>
<ID>IN_0</ID>1431 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k2</lparam></gate>
<gate>
<ID>1238</ID>
<type>DE_TO</type>
<position>628,1491</position>
<input>
<ID>IN_0</ID>1432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID k0</lparam></gate>
<gate>
<ID>1239</ID>
<type>DE_TO</type>
<position>542,1475</position>
<input>
<ID>IN_0</ID>1363 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Subt X</lparam></gate>
<gate>
<ID>1240</ID>
<type>DE_TO</type>
<position>543,1495.5</position>
<input>
<ID>IN_0</ID>1372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AddI X</lparam></gate>
<gate>
<ID>1241</ID>
<type>DE_TO</type>
<position>542,1481</position>
<input>
<ID>IN_0</ID>1351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Output</lparam></gate>
<gate>
<ID>1242</ID>
<type>DE_TO</type>
<position>542,1484</position>
<input>
<ID>IN_0</ID>1352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Halt</lparam></gate>
<gate>
<ID>1243</ID>
<type>DE_TO</type>
<position>541,1490.5</position>
<input>
<ID>IN_0</ID>1338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond1</lparam></gate>
<gate>
<ID>1244</ID>
<type>DA_FROM</type>
<position>701.5,1488</position>
<input>
<ID>IN_0</ID>1346 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1245</ID>
<type>DA_FROM</type>
<position>701.5,1486</position>
<input>
<ID>IN_0</ID>1348 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1246</ID>
<type>DA_FROM</type>
<position>701.5,1484</position>
<input>
<ID>IN_0</ID>1350 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1247</ID>
<type>DA_FROM</type>
<position>701.5,1482</position>
<input>
<ID>IN_0</ID>1362 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1248</ID>
<type>DA_FROM</type>
<position>693,1497</position>
<input>
<ID>IN_0</ID>1364 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1249</ID>
<type>DE_TO</type>
<position>541,1493</position>
<input>
<ID>IN_0</ID>1358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Jump X</lparam></gate>
<gate>
<ID>1250</ID>
<type>AA_TOGGLE</type>
<position>513.5,1481</position>
<output>
<ID>OUT_0</ID>1353 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1251</ID>
<type>DA_FROM</type>
<position>512,1472</position>
<input>
<ID>IN_0</ID>1354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC3</lparam></gate>
<gate>
<ID>1252</ID>
<type>DA_FROM</type>
<position>688,1434</position>
<input>
<ID>IN_0</ID>1359 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MemR</lparam></gate>
<gate>
<ID>1253</ID>
<type>DA_FROM</type>
<position>512,1469</position>
<input>
<ID>IN_0</ID>1355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC2</lparam></gate>
<gate>
<ID>1254</ID>
<type>DA_FROM</type>
<position>512,1466</position>
<input>
<ID>IN_0</ID>1356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC1</lparam></gate>
<gate>
<ID>1255</ID>
<type>DA_FROM</type>
<position>512,1463</position>
<input>
<ID>IN_0</ID>1357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC0</lparam></gate>
<gate>
<ID>1256</ID>
<type>DA_FROM</type>
<position>693,1495</position>
<input>
<ID>IN_0</ID>1365 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1257</ID>
<type>DA_FROM</type>
<position>693,1493</position>
<input>
<ID>IN_0</ID>1366 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1258</ID>
<type>DA_FROM</type>
<position>693,1491</position>
<input>
<ID>IN_0</ID>1367 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1259</ID>
<type>DA_FROM</type>
<position>693,1489</position>
<input>
<ID>IN_0</ID>1368 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1260</ID>
<type>DA_FROM</type>
<position>687.5,1430</position>
<input>
<ID>IN_0</ID>1616 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MemClk</lparam></gate>
<gate>
<ID>1261</ID>
<type>AM_REGISTER16</type>
<position>595.5,1449.5</position>
<input>
<ID>IN_0</ID>1762 </input>
<input>
<ID>IN_1</ID>1763 </input>
<input>
<ID>IN_10</ID>1772 </input>
<input>
<ID>IN_11</ID>1773 </input>
<input>
<ID>IN_12</ID>1774 </input>
<input>
<ID>IN_13</ID>1775 </input>
<input>
<ID>IN_14</ID>1776 </input>
<input>
<ID>IN_15</ID>1777 </input>
<input>
<ID>IN_2</ID>1764 </input>
<input>
<ID>IN_3</ID>1765 </input>
<input>
<ID>IN_4</ID>1766 </input>
<input>
<ID>IN_5</ID>1767 </input>
<input>
<ID>IN_6</ID>1768 </input>
<input>
<ID>IN_7</ID>1769 </input>
<input>
<ID>IN_8</ID>1770 </input>
<input>
<ID>IN_9</ID>1771 </input>
<output>
<ID>OUT_0</ID>1432 </output>
<output>
<ID>OUT_1</ID>1424 </output>
<output>
<ID>OUT_10</ID>1427 </output>
<output>
<ID>OUT_11</ID>1420 </output>
<output>
<ID>OUT_12</ID>1426 </output>
<output>
<ID>OUT_13</ID>1419 </output>
<output>
<ID>OUT_14</ID>1425 </output>
<output>
<ID>OUT_15</ID>1418 </output>
<output>
<ID>OUT_2</ID>1431 </output>
<output>
<ID>OUT_3</ID>1423 </output>
<output>
<ID>OUT_4</ID>1430 </output>
<output>
<ID>OUT_5</ID>1422 </output>
<output>
<ID>OUT_6</ID>1429 </output>
<output>
<ID>OUT_7</ID>1421 </output>
<output>
<ID>OUT_8</ID>1428 </output>
<output>
<ID>OUT_9</ID>1417 </output>
<input>
<ID>clear</ID>1451 </input>
<input>
<ID>clock</ID>1450 </input>
<input>
<ID>load</ID>1493 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1262</ID>
<type>DA_FROM</type>
<position>693,1487</position>
<input>
<ID>IN_0</ID>1369 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1263</ID>
<type>AA_LABEL</type>
<position>598,1474.5</position>
<gparam>LABEL_TEXT ACCUMULATOR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>1264</ID>
<type>DA_FROM</type>
<position>693,1485</position>
<input>
<ID>IN_0</ID>1370 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1265</ID>
<type>DA_FROM</type>
<position>693,1483</position>
<input>
<ID>IN_0</ID>1371 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1266</ID>
<type>AA_AND2</type>
<position>566,1513.5</position>
<input>
<ID>IN_0</ID>1374 </input>
<input>
<ID>IN_1</ID>1390 </input>
<output>
<ID>OUT</ID>1393 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1267</ID>
<type>AA_AND2</type>
<position>565.5,1501.5</position>
<input>
<ID>IN_0</ID>1398 </input>
<input>
<ID>IN_1</ID>1397 </input>
<output>
<ID>OUT</ID>1399 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1268</ID>
<type>AE_SMALL_INVERTER</type>
<position>561,1506</position>
<input>
<ID>IN_0</ID>1374 </input>
<output>
<ID>OUT_0</ID>1398 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1269</ID>
<type>AA_TOGGLE</type>
<position>555.5,1514.5</position>
<output>
<ID>OUT_0</ID>1374 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1270</ID>
<type>AE_OR2</type>
<position>574,1505.5</position>
<input>
<ID>IN_0</ID>1393 </input>
<input>
<ID>IN_1</ID>1399 </input>
<output>
<ID>OUT</ID>1392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1271</ID>
<type>DE_TO</type>
<position>542,1462.5</position>
<input>
<ID>IN_0</ID>1339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JnS</lparam></gate>
<gate>
<ID>1272</ID>
<type>AA_LABEL</type>
<position>538.5,1515.5</position>
<gparam>LABEL_TEXT 1-step/0-countinuos</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1273</ID>
<type>AA_LABEL</type>
<position>543.5,1511</position>
<gparam>LABEL_TEXT STEP BY STEP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1274</ID>
<type>AA_LABEL</type>
<position>548,1506.5</position>
<gparam>LABEL_TEXT RESET</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1275</ID>
<type>DA_FROM</type>
<position>560,1457</position>
<input>
<ID>IN_0</ID>1746 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>1276</ID>
<type>DA_FROM</type>
<position>560,1455</position>
<input>
<ID>IN_0</ID>1747 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>1277</ID>
<type>DA_FROM</type>
<position>560,1453</position>
<input>
<ID>IN_0</ID>1748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>1278</ID>
<type>DA_FROM</type>
<position>560,1451</position>
<input>
<ID>IN_0</ID>1749 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>1279</ID>
<type>DA_FROM</type>
<position>560,1449</position>
<input>
<ID>IN_0</ID>1750 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>1280</ID>
<type>DA_FROM</type>
<position>560,1447</position>
<input>
<ID>IN_0</ID>1751 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>1281</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>686,1489.5</position>
<input>
<ID>ENABLE_0</ID>1378 </input>
<input>
<ID>IN_0</ID>1542 </input>
<input>
<ID>IN_1</ID>1534 </input>
<input>
<ID>IN_10</ID>1537 </input>
<input>
<ID>IN_11</ID>1530 </input>
<input>
<ID>IN_12</ID>1536 </input>
<input>
<ID>IN_13</ID>1529 </input>
<input>
<ID>IN_14</ID>1535 </input>
<input>
<ID>IN_15</ID>1528 </input>
<input>
<ID>IN_2</ID>1541 </input>
<input>
<ID>IN_3</ID>1533 </input>
<input>
<ID>IN_4</ID>1540 </input>
<input>
<ID>IN_5</ID>1532 </input>
<input>
<ID>IN_6</ID>1539 </input>
<input>
<ID>IN_7</ID>1531 </input>
<input>
<ID>IN_8</ID>1538 </input>
<input>
<ID>IN_9</ID>1527 </input>
<output>
<ID>OUT_0</ID>1362 </output>
<output>
<ID>OUT_1</ID>1371 </output>
<output>
<ID>OUT_10</ID>1344 </output>
<output>
<ID>OUT_11</ID>1366 </output>
<output>
<ID>OUT_12</ID>1343 </output>
<output>
<ID>OUT_13</ID>1365 </output>
<output>
<ID>OUT_14</ID>1342 </output>
<output>
<ID>OUT_15</ID>1364 </output>
<output>
<ID>OUT_2</ID>1350 </output>
<output>
<ID>OUT_3</ID>1370 </output>
<output>
<ID>OUT_4</ID>1348 </output>
<output>
<ID>OUT_5</ID>1369 </output>
<output>
<ID>OUT_6</ID>1346 </output>
<output>
<ID>OUT_7</ID>1368 </output>
<output>
<ID>OUT_8</ID>1345 </output>
<output>
<ID>OUT_9</ID>1367 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1282</ID>
<type>DA_FROM</type>
<position>696,1501</position>
<input>
<ID>IN_0</ID>1378 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MDBR</lparam></gate>
<gate>
<ID>1283</ID>
<type>DA_FROM</type>
<position>559.5,1445</position>
<input>
<ID>IN_0</ID>1752 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>1284</ID>
<type>DA_FROM</type>
<position>559,1443</position>
<input>
<ID>IN_0</ID>1753 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>1285</ID>
<type>DA_FROM</type>
<position>551.5,1444</position>
<input>
<ID>IN_0</ID>1756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>1286</ID>
<type>DA_FROM</type>
<position>551.5,1442</position>
<input>
<ID>IN_0</ID>1757 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>1287</ID>
<type>DA_FROM</type>
<position>551.5,1456</position>
<input>
<ID>IN_0</ID>1758 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>1288</ID>
<type>DA_FROM</type>
<position>572,1484</position>
<input>
<ID>IN_0</ID>1341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACW1</lparam></gate>
<gate>
<ID>1289</ID>
<type>DA_FROM</type>
<position>551.5,1454</position>
<input>
<ID>IN_0</ID>1759 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>1290</ID>
<type>DA_FROM</type>
<position>551.5,1452</position>
<input>
<ID>IN_0</ID>1760 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>1291</ID>
<type>AA_TOGGLE</type>
<position>565.5,1463</position>
<output>
<ID>OUT_0</ID>1380 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1292</ID>
<type>AA_TOGGLE</type>
<position>565.5,1465</position>
<output>
<ID>OUT_0</ID>1381 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1293</ID>
<type>AA_TOGGLE</type>
<position>565.5,1467</position>
<output>
<ID>OUT_0</ID>1379 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1294</ID>
<type>AA_TOGGLE</type>
<position>565.5,1469</position>
<output>
<ID>OUT_0</ID>1382 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1295</ID>
<type>AA_TOGGLE</type>
<position>565.5,1471</position>
<output>
<ID>OUT_0</ID>1383 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1296</ID>
<type>AA_TOGGLE</type>
<position>565.5,1473</position>
<output>
<ID>OUT_0</ID>1384 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1297</ID>
<type>AA_TOGGLE</type>
<position>565.5,1475</position>
<output>
<ID>OUT_0</ID>1385 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1298</ID>
<type>AA_TOGGLE</type>
<position>565.5,1477</position>
<output>
<ID>OUT_0</ID>1386 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1299</ID>
<type>AA_TOGGLE</type>
<position>569,1464</position>
<output>
<ID>OUT_0</ID>1387 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1300</ID>
<type>AA_TOGGLE</type>
<position>569,1466</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1301</ID>
<type>AA_TOGGLE</type>
<position>569,1468</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1302</ID>
<type>AA_TOGGLE</type>
<position>569,1470</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1303</ID>
<type>AA_TOGGLE</type>
<position>569,1472</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1304</ID>
<type>AA_TOGGLE</type>
<position>569,1474</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1305</ID>
<type>AA_TOGGLE</type>
<position>569,1476</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1306</ID>
<type>AA_TOGGLE</type>
<position>569,1478</position>
<output>
<ID>OUT_0</ID>1388 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1307</ID>
<type>DA_FROM</type>
<position>551.5,1450</position>
<input>
<ID>IN_0</ID>1761 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>1308</ID>
<type>DA_FROM</type>
<position>651,1489.5</position>
<input>
<ID>IN_0</ID>1375 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALUS</lparam></gate>
<gate>
<ID>1309</ID>
<type>DA_FROM</type>
<position>551.5,1448</position>
<input>
<ID>IN_0</ID>1754 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>1310</ID>
<type>DA_FROM</type>
<position>551.5,1446</position>
<input>
<ID>IN_0</ID>1755 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>1311</ID>
<type>DA_FROM</type>
<position>642.5,1424</position>
<input>
<ID>IN_0</ID>1401 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1312</ID>
<type>DE_TO</type>
<position>634,1483</position>
<input>
<ID>IN_0</ID>1321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC15</lparam></gate>
<gate>
<ID>1313</ID>
<type>DE_TO</type>
<position>634,1481</position>
<input>
<ID>IN_0</ID>1322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC13</lparam></gate>
<gate>
<ID>1314</ID>
<type>DE_TO</type>
<position>634,1479</position>
<input>
<ID>IN_0</ID>1323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC11</lparam></gate>
<gate>
<ID>1315</ID>
<type>DE_TO</type>
<position>634,1477</position>
<input>
<ID>IN_0</ID>1324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC9</lparam></gate>
<gate>
<ID>1316</ID>
<type>DE_TO</type>
<position>634,1475</position>
<input>
<ID>IN_0</ID>1325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC7</lparam></gate>
<gate>
<ID>1317</ID>
<type>DE_TO</type>
<position>634,1473</position>
<input>
<ID>IN_0</ID>1326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC5</lparam></gate>
<gate>
<ID>1318</ID>
<type>DE_TO</type>
<position>634,1471</position>
<input>
<ID>IN_0</ID>1327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC3</lparam></gate>
<gate>
<ID>1319</ID>
<type>DE_TO</type>
<position>634,1469</position>
<input>
<ID>IN_0</ID>1328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC1</lparam></gate>
<gate>
<ID>1320</ID>
<type>DE_TO</type>
<position>627,1482</position>
<input>
<ID>IN_0</ID>1329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC14</lparam></gate>
<gate>
<ID>1321</ID>
<type>DE_TO</type>
<position>627,1480</position>
<input>
<ID>IN_0</ID>1330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC12</lparam></gate>
<gate>
<ID>1322</ID>
<type>DE_TO</type>
<position>627,1478</position>
<input>
<ID>IN_0</ID>1331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC10</lparam></gate>
<gate>
<ID>1323</ID>
<type>DE_TO</type>
<position>627,1476</position>
<input>
<ID>IN_0</ID>1332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC8</lparam></gate>
<gate>
<ID>1324</ID>
<type>DE_TO</type>
<position>627,1474</position>
<input>
<ID>IN_0</ID>1333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC6</lparam></gate>
<gate>
<ID>1325</ID>
<type>DE_TO</type>
<position>627,1472</position>
<input>
<ID>IN_0</ID>1334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC4</lparam></gate>
<gate>
<ID>1326</ID>
<type>DE_TO</type>
<position>627,1470</position>
<input>
<ID>IN_0</ID>1335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC2</lparam></gate>
<gate>
<ID>1327</ID>
<type>DE_TO</type>
<position>627,1468</position>
<input>
<ID>IN_0</ID>1336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC0</lparam></gate>
<gate>
<ID>1328</ID>
<type>DA_FROM</type>
<position>642.5,1422</position>
<input>
<ID>IN_0</ID>1400 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1329</ID>
<type>DA_FROM</type>
<position>636,1423</position>
<input>
<ID>IN_0</ID>1408 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1330</ID>
<type>DA_FROM</type>
<position>636,1421</position>
<input>
<ID>IN_0</ID>1409 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1331</ID>
<type>DA_FROM</type>
<position>636,1435</position>
<input>
<ID>IN_0</ID>1410 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1332</ID>
<type>DA_FROM</type>
<position>636,1433</position>
<input>
<ID>IN_0</ID>1411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1333</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>621,1449.5</position>
<input>
<ID>ENABLE_0</ID>1433 </input>
<input>
<ID>IN_0</ID>1432 </input>
<input>
<ID>IN_1</ID>1424 </input>
<input>
<ID>IN_10</ID>1427 </input>
<input>
<ID>IN_11</ID>1420 </input>
<input>
<ID>IN_12</ID>1426 </input>
<input>
<ID>IN_13</ID>1419 </input>
<input>
<ID>IN_14</ID>1425 </input>
<input>
<ID>IN_15</ID>1418 </input>
<input>
<ID>IN_2</ID>1431 </input>
<input>
<ID>IN_3</ID>1423 </input>
<input>
<ID>IN_4</ID>1430 </input>
<input>
<ID>IN_5</ID>1422 </input>
<input>
<ID>IN_6</ID>1429 </input>
<input>
<ID>IN_7</ID>1421 </input>
<input>
<ID>IN_8</ID>1428 </input>
<input>
<ID>IN_9</ID>1417 </input>
<output>
<ID>OUT_0</ID>1441 </output>
<output>
<ID>OUT_1</ID>1444 </output>
<output>
<ID>OUT_10</ID>1436 </output>
<output>
<ID>OUT_11</ID>1447 </output>
<output>
<ID>OUT_12</ID>1435 </output>
<output>
<ID>OUT_13</ID>1448 </output>
<output>
<ID>OUT_14</ID>1434 </output>
<output>
<ID>OUT_15</ID>1449 </output>
<output>
<ID>OUT_2</ID>1440 </output>
<output>
<ID>OUT_3</ID>1443 </output>
<output>
<ID>OUT_4</ID>1439 </output>
<output>
<ID>OUT_5</ID>1442 </output>
<output>
<ID>OUT_6</ID>1438 </output>
<output>
<ID>OUT_7</ID>1445 </output>
<output>
<ID>OUT_8</ID>1437 </output>
<output>
<ID>OUT_9</ID>1446 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1334</ID>
<type>DA_FROM</type>
<position>636,1431</position>
<input>
<ID>IN_0</ID>1412 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1335</ID>
<type>DA_FROM</type>
<position>621,1462</position>
<input>
<ID>IN_0</ID>1433 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID ACS</lparam></gate>
<gate>
<ID>1336</ID>
<type>DE_TO</type>
<position>634.5,1457</position>
<input>
<ID>IN_0</ID>1449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1337</ID>
<type>DE_TO</type>
<position>634.5,1455</position>
<input>
<ID>IN_0</ID>1448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1338</ID>
<type>DE_TO</type>
<position>634.5,1453</position>
<input>
<ID>IN_0</ID>1447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1339</ID>
<type>DE_TO</type>
<position>634.5,1451</position>
<input>
<ID>IN_0</ID>1446 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1340</ID>
<type>DE_TO</type>
<position>634.5,1449</position>
<input>
<ID>IN_0</ID>1445 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1341</ID>
<type>DE_TO</type>
<position>634.5,1447</position>
<input>
<ID>IN_0</ID>1442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1342</ID>
<type>DE_TO</type>
<position>634.5,1445</position>
<input>
<ID>IN_0</ID>1443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1343</ID>
<type>DE_TO</type>
<position>634.5,1443</position>
<input>
<ID>IN_0</ID>1444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1344</ID>
<type>DE_TO</type>
<position>627.5,1456</position>
<input>
<ID>IN_0</ID>1434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1345</ID>
<type>DE_TO</type>
<position>627.5,1454</position>
<input>
<ID>IN_0</ID>1435 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1346</ID>
<type>DE_TO</type>
<position>627.5,1452</position>
<input>
<ID>IN_0</ID>1436 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1347</ID>
<type>DE_TO</type>
<position>627.5,1450</position>
<input>
<ID>IN_0</ID>1437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1348</ID>
<type>DE_TO</type>
<position>627.5,1448</position>
<input>
<ID>IN_0</ID>1438 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1349</ID>
<type>DE_TO</type>
<position>627.5,1446</position>
<input>
<ID>IN_0</ID>1439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1350</ID>
<type>DE_TO</type>
<position>627.5,1444</position>
<input>
<ID>IN_0</ID>1440 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1351</ID>
<type>DE_TO</type>
<position>627.5,1442</position>
<input>
<ID>IN_0</ID>1441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1352</ID>
<type>DA_FROM</type>
<position>636,1429</position>
<input>
<ID>IN_0</ID>1413 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1353</ID>
<type>DA_FROM</type>
<position>636,1427</position>
<input>
<ID>IN_0</ID>1414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1354</ID>
<type>AE_OR2</type>
<position>589.5,1437</position>
<input>
<ID>IN_0</ID>1452 </input>
<input>
<ID>IN_1</ID>1453 </input>
<output>
<ID>OUT</ID>1450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1355</ID>
<type>DA_FROM</type>
<position>636,1425</position>
<input>
<ID>IN_0</ID>1415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1356</ID>
<type>AE_OR2</type>
<position>605,1437</position>
<input>
<ID>IN_0</ID>1455 </input>
<input>
<ID>IN_1</ID>1454 </input>
<output>
<ID>OUT</ID>1451 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1357</ID>
<type>DA_FROM</type>
<position>642.5,1436</position>
<input>
<ID>IN_0</ID>1402 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1358</ID>
<type>DA_FROM</type>
<position>579.5,1438</position>
<input>
<ID>IN_0</ID>1452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACW</lparam></gate>
<gate>
<ID>1359</ID>
<type>DA_FROM</type>
<position>642.5,1434</position>
<input>
<ID>IN_0</ID>1403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1360</ID>
<type>DA_FROM</type>
<position>576,1436</position>
<input>
<ID>IN_0</ID>1453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1361</ID>
<type>DA_FROM</type>
<position>642.5,1432</position>
<input>
<ID>IN_0</ID>1404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1362</ID>
<type>DA_FROM</type>
<position>615.5,1438</position>
<input>
<ID>IN_0</ID>1454 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ACS</lparam></gate>
<gate>
<ID>1363</ID>
<type>DA_FROM</type>
<position>642.5,1430</position>
<input>
<ID>IN_0</ID>1405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1364</ID>
<type>DA_FROM</type>
<position>642.5,1428</position>
<input>
<ID>IN_0</ID>1406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1365</ID>
<type>DA_FROM</type>
<position>642.5,1426</position>
<input>
<ID>IN_0</ID>1407 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1366</ID>
<type>AA_LABEL</type>
<position>605.5,1427</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1367</ID>
<type>AA_LABEL</type>
<position>665.5,1448</position>
<gparam>LABEL_TEXT Memory Adres Register     Memory</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1368</ID>
<type>DA_FROM</type>
<position>590.5,1402</position>
<input>
<ID>IN_0</ID>1462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1369</ID>
<type>DA_FROM</type>
<position>590.5,1400</position>
<input>
<ID>IN_0</ID>1461 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1370</ID>
<type>DA_FROM</type>
<position>582,1401</position>
<input>
<ID>IN_0</ID>1469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1371</ID>
<type>DA_FROM</type>
<position>582,1399</position>
<input>
<ID>IN_0</ID>1468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1372</ID>
<type>DA_FROM</type>
<position>582,1413</position>
<input>
<ID>IN_0</ID>1467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1373</ID>
<type>DA_FROM</type>
<position>582,1411</position>
<input>
<ID>IN_0</ID>1466 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1374</ID>
<type>DA_FROM</type>
<position>582,1409</position>
<input>
<ID>IN_0</ID>1470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1375</ID>
<type>DA_FROM</type>
<position>582,1407</position>
<input>
<ID>IN_0</ID>1465 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1376</ID>
<type>DA_FROM</type>
<position>582,1405</position>
<input>
<ID>IN_0</ID>1464 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1377</ID>
<type>DA_FROM</type>
<position>610,1436</position>
<input>
<ID>IN_0</ID>1455 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1378</ID>
<type>DA_FROM</type>
<position>582,1403</position>
<input>
<ID>IN_0</ID>1463 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1379</ID>
<type>DA_FROM</type>
<position>590.5,1414</position>
<input>
<ID>IN_0</ID>1460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1380</ID>
<type>DA_FROM</type>
<position>590.5,1412</position>
<input>
<ID>IN_0</ID>1459 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1381</ID>
<type>DA_FROM</type>
<position>590.5,1410</position>
<input>
<ID>IN_0</ID>1458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1382</ID>
<type>DA_FROM</type>
<position>590.5,1408</position>
<input>
<ID>IN_0</ID>1457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1383</ID>
<type>DA_FROM</type>
<position>590.5,1406</position>
<input>
<ID>IN_0</ID>1456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1384</ID>
<type>DA_FROM</type>
<position>590.5,1404</position>
<input>
<ID>IN_0</ID>1416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1385</ID>
<type>DE_TO</type>
<position>621,1414</position>
<input>
<ID>IN_0</ID>1483 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1386</ID>
<type>DE_TO</type>
<position>621,1412</position>
<input>
<ID>IN_0</ID>1482 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1387</ID>
<type>DE_TO</type>
<position>621,1410</position>
<input>
<ID>IN_0</ID>1481 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1388</ID>
<type>DE_TO</type>
<position>621,1408</position>
<input>
<ID>IN_0</ID>1480 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1389</ID>
<type>DE_TO</type>
<position>621,1406</position>
<input>
<ID>IN_0</ID>1479 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1390</ID>
<type>DE_TO</type>
<position>621,1404</position>
<input>
<ID>IN_0</ID>1484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1391</ID>
<type>DE_TO</type>
<position>621,1402</position>
<input>
<ID>IN_0</ID>1485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1392</ID>
<type>DE_TO</type>
<position>621,1400</position>
<input>
<ID>IN_0</ID>1486 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1393</ID>
<type>DE_TO</type>
<position>613.5,1413</position>
<input>
<ID>IN_0</ID>1472 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1394</ID>
<type>DE_TO</type>
<position>613.5,1411</position>
<input>
<ID>IN_0</ID>1471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1395</ID>
<type>DE_TO</type>
<position>613.5,1409</position>
<input>
<ID>IN_0</ID>1478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1396</ID>
<type>DE_TO</type>
<position>613.5,1407</position>
<input>
<ID>IN_0</ID>1477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1397</ID>
<type>DE_TO</type>
<position>613.5,1405</position>
<input>
<ID>IN_0</ID>1476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1398</ID>
<type>DE_TO</type>
<position>613.5,1403</position>
<input>
<ID>IN_0</ID>1475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1399</ID>
<type>DE_TO</type>
<position>613.5,1401</position>
<input>
<ID>IN_0</ID>1474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1400</ID>
<type>DE_TO</type>
<position>613.5,1399</position>
<input>
<ID>IN_0</ID>1473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1401</ID>
<type>DA_FROM</type>
<position>587,1422.5</position>
<input>
<ID>IN_0</ID>1488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCL</lparam></gate>
<gate>
<ID>1402</ID>
<type>AE_SMALL_INVERTER</type>
<position>599,1419.5</position>
<input>
<ID>IN_0</ID>1488 </input>
<output>
<ID>OUT_0</ID>1487 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1403</ID>
<type>EE_VDD</type>
<position>600,1422.5</position>
<output>
<ID>OUT_0</ID>1489 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1404</ID>
<type>FF_GND</type>
<position>602,1422.5</position>
<output>
<ID>OUT_0</ID>1490 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1405</ID>
<type>EE_VDD</type>
<position>649.5,1441.5</position>
<output>
<ID>OUT_0</ID>1491 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1406</ID>
<type>EE_VDD</type>
<position>667,1482.5</position>
<output>
<ID>OUT_0</ID>1492 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1407</ID>
<type>EE_VDD</type>
<position>594.5,1463.5</position>
<output>
<ID>OUT_0</ID>1493 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1408</ID>
<type>DA_FROM</type>
<position>714,1473.5</position>
<input>
<ID>IN_0</ID>1509 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1409</ID>
<type>DA_FROM</type>
<position>714,1471.5</position>
<input>
<ID>IN_0</ID>1504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1410</ID>
<type>DA_FROM</type>
<position>714,1469.5</position>
<input>
<ID>IN_0</ID>1503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1411</ID>
<type>DA_FROM</type>
<position>714,1467.5</position>
<input>
<ID>IN_0</ID>1502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1412</ID>
<type>DA_FROM</type>
<position>722.5,1478.5</position>
<input>
<ID>IN_0</ID>1499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1413</ID>
<type>DA_FROM</type>
<position>722.5,1476.5</position>
<input>
<ID>IN_0</ID>1498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1414</ID>
<type>DA_FROM</type>
<position>722.5,1474.5</position>
<input>
<ID>IN_0</ID>1497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1415</ID>
<type>DA_FROM</type>
<position>722.5,1472.5</position>
<input>
<ID>IN_0</ID>1496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1416</ID>
<type>DA_FROM</type>
<position>722.5,1470.5</position>
<input>
<ID>IN_0</ID>1495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1417</ID>
<type>DA_FROM</type>
<position>722.5,1468.5</position>
<input>
<ID>IN_0</ID>1494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1418</ID>
<type>DE_TO</type>
<position>757.5,1478.5</position>
<input>
<ID>IN_0</ID>1554 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1419</ID>
<type>DE_TO</type>
<position>757.5,1476.5</position>
<input>
<ID>IN_0</ID>1553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1420</ID>
<type>DE_TO</type>
<position>757.5,1474.5</position>
<input>
<ID>IN_0</ID>1552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1421</ID>
<type>DE_TO</type>
<position>757.5,1472.5</position>
<input>
<ID>IN_0</ID>1551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1422</ID>
<type>DE_TO</type>
<position>757.5,1470.5</position>
<input>
<ID>IN_0</ID>1550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1423</ID>
<type>DE_TO</type>
<position>757.5,1468.5</position>
<input>
<ID>IN_0</ID>1555 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1424</ID>
<type>DE_TO</type>
<position>757.5,1466.5</position>
<input>
<ID>IN_0</ID>1556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1425</ID>
<type>DE_TO</type>
<position>757.5,1464.5</position>
<input>
<ID>IN_0</ID>1557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1426</ID>
<type>DE_TO</type>
<position>750,1477.5</position>
<input>
<ID>IN_0</ID>1543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1427</ID>
<type>DE_TO</type>
<position>750,1475.5</position>
<input>
<ID>IN_0</ID>1510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1428</ID>
<type>DE_TO</type>
<position>750,1473.5</position>
<input>
<ID>IN_0</ID>1549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1429</ID>
<type>DE_TO</type>
<position>750,1471.5</position>
<input>
<ID>IN_0</ID>1548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1430</ID>
<type>DE_TO</type>
<position>750,1469.5</position>
<input>
<ID>IN_0</ID>1547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1431</ID>
<type>DA_FROM</type>
<position>660,1466.5</position>
<input>
<ID>IN_0</ID>1517 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1432</ID>
<type>DA_FROM</type>
<position>660,1464.5</position>
<input>
<ID>IN_0</ID>1518 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1433</ID>
<type>DA_FROM</type>
<position>653.5,1465.5</position>
<input>
<ID>IN_0</ID>1519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1434</ID>
<type>DA_FROM</type>
<position>653.5,1463.5</position>
<input>
<ID>IN_0</ID>1520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1435</ID>
<type>DA_FROM</type>
<position>653.5,1477.5</position>
<input>
<ID>IN_0</ID>1521 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1436</ID>
<type>DA_FROM</type>
<position>672.5,1457.5</position>
<input>
<ID>IN_0</ID>1561 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1437</ID>
<type>DA_FROM</type>
<position>653.5,1475.5</position>
<input>
<ID>IN_0</ID>1522 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1438</ID>
<type>DA_FROM</type>
<position>653.5,1473.5</position>
<input>
<ID>IN_0</ID>1523 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D10</lparam></gate>
<gate>
<ID>1439</ID>
<type>DA_FROM</type>
<position>653.5,1471.5</position>
<input>
<ID>IN_0</ID>1524 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D8</lparam></gate>
<gate>
<ID>1440</ID>
<type>DA_FROM</type>
<position>653.5,1469.5</position>
<input>
<ID>IN_0</ID>1525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>1441</ID>
<type>DA_FROM</type>
<position>653.5,1467.5</position>
<input>
<ID>IN_0</ID>1526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1442</ID>
<type>DE_TO</type>
<position>698.5,1478.5</position>
<input>
<ID>IN_0</ID>1528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR15</lparam></gate>
<gate>
<ID>1443</ID>
<type>DE_TO</type>
<position>698.5,1476.5</position>
<input>
<ID>IN_0</ID>1529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR13</lparam></gate>
<gate>
<ID>1444</ID>
<type>DE_TO</type>
<position>698.5,1474.5</position>
<input>
<ID>IN_0</ID>1530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR11</lparam></gate>
<gate>
<ID>1445</ID>
<type>DE_TO</type>
<position>698.5,1472.5</position>
<input>
<ID>IN_0</ID>1527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR9</lparam></gate>
<gate>
<ID>1446</ID>
<type>DE_TO</type>
<position>698.5,1470.5</position>
<input>
<ID>IN_0</ID>1531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR7</lparam></gate>
<gate>
<ID>1447</ID>
<type>DE_TO</type>
<position>698.5,1468.5</position>
<input>
<ID>IN_0</ID>1532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR5</lparam></gate>
<gate>
<ID>1448</ID>
<type>DE_TO</type>
<position>698.5,1466.5</position>
<input>
<ID>IN_0</ID>1533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR3</lparam></gate>
<gate>
<ID>1449</ID>
<type>DE_TO</type>
<position>698.5,1464.5</position>
<input>
<ID>IN_0</ID>1534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR1</lparam></gate>
<gate>
<ID>1450</ID>
<type>DE_TO</type>
<position>687,1477.5</position>
<input>
<ID>IN_0</ID>1535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR14</lparam></gate>
<gate>
<ID>1451</ID>
<type>DE_TO</type>
<position>687,1475.5</position>
<input>
<ID>IN_0</ID>1536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR12</lparam></gate>
<gate>
<ID>1452</ID>
<type>DE_TO</type>
<position>687,1473.5</position>
<input>
<ID>IN_0</ID>1537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR10</lparam></gate>
<gate>
<ID>1453</ID>
<type>DE_TO</type>
<position>687,1471.5</position>
<input>
<ID>IN_0</ID>1538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR8</lparam></gate>
<gate>
<ID>1454</ID>
<type>DE_TO</type>
<position>687,1469.5</position>
<input>
<ID>IN_0</ID>1539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR6</lparam></gate>
<gate>
<ID>1455</ID>
<type>DE_TO</type>
<position>687,1467.5</position>
<input>
<ID>IN_0</ID>1540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR4</lparam></gate>
<gate>
<ID>1456</ID>
<type>DE_TO</type>
<position>687,1465.5</position>
<input>
<ID>IN_0</ID>1541 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR2</lparam></gate>
<gate>
<ID>1457</ID>
<type>DE_TO</type>
<position>687,1463.5</position>
<input>
<ID>IN_0</ID>1542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR0</lparam></gate>
<gate>
<ID>1458</ID>
<type>AM_REGISTER16</type>
<position>668,1471</position>
<input>
<ID>IN_0</ID>1520 </input>
<input>
<ID>IN_1</ID>1518 </input>
<input>
<ID>IN_10</ID>1523 </input>
<input>
<ID>IN_11</ID>1513 </input>
<input>
<ID>IN_12</ID>1522 </input>
<input>
<ID>IN_13</ID>1512 </input>
<input>
<ID>IN_14</ID>1521 </input>
<input>
<ID>IN_15</ID>1511 </input>
<input>
<ID>IN_2</ID>1519 </input>
<input>
<ID>IN_3</ID>1517 </input>
<input>
<ID>IN_4</ID>1526 </input>
<input>
<ID>IN_5</ID>1516 </input>
<input>
<ID>IN_6</ID>1525 </input>
<input>
<ID>IN_7</ID>1515 </input>
<input>
<ID>IN_8</ID>1524 </input>
<input>
<ID>IN_9</ID>1514 </input>
<output>
<ID>OUT_0</ID>1542 </output>
<output>
<ID>OUT_1</ID>1534 </output>
<output>
<ID>OUT_10</ID>1537 </output>
<output>
<ID>OUT_11</ID>1530 </output>
<output>
<ID>OUT_12</ID>1536 </output>
<output>
<ID>OUT_13</ID>1529 </output>
<output>
<ID>OUT_14</ID>1535 </output>
<output>
<ID>OUT_15</ID>1528 </output>
<output>
<ID>OUT_2</ID>1541 </output>
<output>
<ID>OUT_3</ID>1533 </output>
<output>
<ID>OUT_4</ID>1540 </output>
<output>
<ID>OUT_5</ID>1532 </output>
<output>
<ID>OUT_6</ID>1539 </output>
<output>
<ID>OUT_7</ID>1531 </output>
<output>
<ID>OUT_8</ID>1538 </output>
<output>
<ID>OUT_9</ID>1527 </output>
<input>
<ID>clear</ID>1561 </input>
<input>
<ID>clock</ID>1558 </input>
<input>
<ID>load</ID>1492 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1459</ID>
<type>DE_TO</type>
<position>750,1467.5</position>
<input>
<ID>IN_0</ID>1546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>1460</ID>
<type>DE_TO</type>
<position>750,1465.5</position>
<input>
<ID>IN_0</ID>1545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1461</ID>
<type>DE_TO</type>
<position>750,1463.5</position>
<input>
<ID>IN_0</ID>1544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1462</ID>
<type>DA_FROM</type>
<position>734,1456.5</position>
<input>
<ID>IN_0</ID>1606 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1463</ID>
<type>AM_REGISTER16</type>
<position>731,1471</position>
<input>
<ID>IN_0</ID>1507 </input>
<input>
<ID>IN_1</ID>1500 </input>
<input>
<ID>IN_10</ID>1509 </input>
<input>
<ID>IN_11</ID>1497 </input>
<input>
<ID>IN_12</ID>1505 </input>
<input>
<ID>IN_13</ID>1498 </input>
<input>
<ID>IN_14</ID>1506 </input>
<input>
<ID>IN_15</ID>1499 </input>
<input>
<ID>IN_2</ID>1508 </input>
<input>
<ID>IN_3</ID>1501 </input>
<input>
<ID>IN_4</ID>1502 </input>
<input>
<ID>IN_5</ID>1494 </input>
<input>
<ID>IN_6</ID>1503 </input>
<input>
<ID>IN_7</ID>1495 </input>
<input>
<ID>IN_8</ID>1504 </input>
<input>
<ID>IN_9</ID>1496 </input>
<output>
<ID>OUT_0</ID>1586 </output>
<output>
<ID>OUT_1</ID>1580 </output>
<output>
<ID>OUT_10</ID>1581 </output>
<output>
<ID>OUT_11</ID>1576 </output>
<output>
<ID>OUT_12</ID>1609 </output>
<output>
<ID>OUT_13</ID>1610 </output>
<output>
<ID>OUT_14</ID>1611 </output>
<output>
<ID>OUT_15</ID>1612 </output>
<output>
<ID>OUT_2</ID>1585 </output>
<output>
<ID>OUT_3</ID>1579 </output>
<output>
<ID>OUT_4</ID>1584 </output>
<output>
<ID>OUT_5</ID>1578 </output>
<output>
<ID>OUT_6</ID>1583 </output>
<output>
<ID>OUT_7</ID>1577 </output>
<output>
<ID>OUT_8</ID>1582 </output>
<output>
<ID>OUT_9</ID>1575 </output>
<input>
<ID>clear</ID>1606 </input>
<input>
<ID>clock</ID>1604 </input>
<input>
<ID>load</ID>1608 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1464</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>743.5,1471</position>
<input>
<ID>ENABLE_0</ID>1607 </input>
<input>
<ID>IN_0</ID>1586 </input>
<input>
<ID>IN_1</ID>1580 </input>
<input>
<ID>IN_10</ID>1581 </input>
<input>
<ID>IN_11</ID>1576 </input>
<input>
<ID>IN_12</ID>1615 </input>
<input>
<ID>IN_13</ID>1615 </input>
<input>
<ID>IN_14</ID>1615 </input>
<input>
<ID>IN_15</ID>1615 </input>
<input>
<ID>IN_2</ID>1585 </input>
<input>
<ID>IN_3</ID>1579 </input>
<input>
<ID>IN_4</ID>1584 </input>
<input>
<ID>IN_5</ID>1578 </input>
<input>
<ID>IN_6</ID>1583 </input>
<input>
<ID>IN_7</ID>1577 </input>
<input>
<ID>IN_8</ID>1582 </input>
<input>
<ID>IN_9</ID>1575 </input>
<output>
<ID>OUT_0</ID>1544 </output>
<output>
<ID>OUT_1</ID>1557 </output>
<output>
<ID>OUT_10</ID>1549 </output>
<output>
<ID>OUT_11</ID>1552 </output>
<output>
<ID>OUT_12</ID>1510 </output>
<output>
<ID>OUT_13</ID>1553 </output>
<output>
<ID>OUT_14</ID>1543 </output>
<output>
<ID>OUT_15</ID>1554 </output>
<output>
<ID>OUT_2</ID>1545 </output>
<output>
<ID>OUT_3</ID>1556 </output>
<output>
<ID>OUT_4</ID>1546 </output>
<output>
<ID>OUT_5</ID>1555 </output>
<output>
<ID>OUT_6</ID>1547 </output>
<output>
<ID>OUT_7</ID>1550 </output>
<output>
<ID>OUT_8</ID>1548 </output>
<output>
<ID>OUT_9</ID>1551 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1465</ID>
<type>DA_FROM</type>
<position>749,1481.5</position>
<input>
<ID>IN_0</ID>1607 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IRS</lparam></gate>
<gate>
<ID>1466</ID>
<type>AE_OR2</type>
<position>726,1456.5</position>
<input>
<ID>IN_0</ID>1613 </input>
<input>
<ID>IN_1</ID>1605 </input>
<output>
<ID>OUT</ID>1604 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1467</ID>
<type>DA_FROM</type>
<position>720,1455.5</position>
<input>
<ID>IN_0</ID>1605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1468</ID>
<type>AE_OR2</type>
<position>662.5,1457.5</position>
<input>
<ID>IN_0</ID>1559 </input>
<input>
<ID>IN_1</ID>1560 </input>
<output>
<ID>OUT</ID>1558 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1469</ID>
<type>DA_FROM</type>
<position>660,1478.5</position>
<input>
<ID>IN_0</ID>1511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D15</lparam></gate>
<gate>
<ID>1470</ID>
<type>DA_FROM</type>
<position>718,1457.5</position>
<input>
<ID>IN_0</ID>1613 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRW</lparam></gate>
<gate>
<ID>1471</ID>
<type>DA_FROM</type>
<position>660,1476.5</position>
<input>
<ID>IN_0</ID>1512 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D13</lparam></gate>
<gate>
<ID>1472</ID>
<type>DA_FROM</type>
<position>660,1474.5</position>
<input>
<ID>IN_0</ID>1513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D11</lparam></gate>
<gate>
<ID>1473</ID>
<type>DA_FROM</type>
<position>654.5,1458.5</position>
<input>
<ID>IN_0</ID>1559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDBW</lparam></gate>
<gate>
<ID>1474</ID>
<type>DA_FROM</type>
<position>660,1472.5</position>
<input>
<ID>IN_0</ID>1514 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D9</lparam></gate>
<gate>
<ID>1475</ID>
<type>DA_FROM</type>
<position>660,1470.5</position>
<input>
<ID>IN_0</ID>1515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>1476</ID>
<type>DA_FROM</type>
<position>660,1468.5</position>
<input>
<ID>IN_0</ID>1516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>1477</ID>
<type>DA_FROM</type>
<position>654.5,1456.5</position>
<input>
<ID>IN_0</ID>1560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1478</ID>
<type>AA_LABEL</type>
<position>721,1488</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1479</ID>
<type>DA_FROM</type>
<position>722.5,1466.5</position>
<input>
<ID>IN_0</ID>1501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1480</ID>
<type>AA_LABEL</type>
<position>688.5,1505</position>
<gparam>LABEL_TEXT MEMORY DATA BUFFER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1481</ID>
<type>DA_FROM</type>
<position>722.5,1464.5</position>
<input>
<ID>IN_0</ID>1500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1482</ID>
<type>AA_TOGGLE</type>
<position>528.5,1407</position>
<output>
<ID>OUT_0</ID>1562 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1483</ID>
<type>DA_FROM</type>
<position>714,1465.5</position>
<input>
<ID>IN_0</ID>1508 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1484</ID>
<type>CC_PULSE</type>
<position>555.5,1506</position>
<output>
<ID>OUT_0</ID>1742 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1485</ID>
<type>DA_FROM</type>
<position>714,1463.5</position>
<input>
<ID>IN_0</ID>1507 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>1486</ID>
<type>DA_FROM</type>
<position>714,1477.5</position>
<input>
<ID>IN_0</ID>1506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D14</lparam></gate>
<gate>
<ID>1487</ID>
<type>DA_FROM</type>
<position>714,1475.5</position>
<input>
<ID>IN_0</ID>1505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D12</lparam></gate>
<gate>
<ID>1488</ID>
<type>EE_VDD</type>
<position>730,1483.5</position>
<output>
<ID>OUT_0</ID>1608 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1489</ID>
<type>DE_TO</type>
<position>538.5,1407</position>
<input>
<ID>IN_0</ID>1562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Start</lparam></gate>
<gate>
<ID>1490</ID>
<type>DE_TO</type>
<position>579,1497</position>
<input>
<ID>IN_0</ID>1742 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>1491</ID>
<type>AE_DFF_LOW</type>
<position>641,1388</position>
<input>
<ID>IN_0</ID>1563 </input>
<output>
<ID>OUTINV_0</ID>1563 </output>
<output>
<ID>OUT_0</ID>1567 </output>
<input>
<ID>clock</ID>1571 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1492</ID>
<type>DE_TO</type>
<position>746.5,1483.5</position>
<input>
<ID>IN_0</ID>1609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC0</lparam></gate>
<gate>
<ID>1493</ID>
<type>DA_FROM</type>
<position>617,1388</position>
<input>
<ID>IN_0</ID>1564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Reset</lparam></gate>
<gate>
<ID>1494</ID>
<type>DE_TO</type>
<position>746.5,1485.5</position>
<input>
<ID>IN_0</ID>1610 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC1</lparam></gate>
<gate>
<ID>1495</ID>
<type>AE_SMALL_INVERTER</type>
<position>623.5,1391</position>
<input>
<ID>IN_0</ID>1564 </input>
<output>
<ID>OUT_0</ID>1565 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1496</ID>
<type>AE_SMALL_INVERTER</type>
<position>628.5,1391</position>
<input>
<ID>IN_0</ID>1565 </input>
<output>
<ID>OUT_0</ID>1566 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1497</ID>
<type>DE_TO</type>
<position>746.5,1487.5</position>
<input>
<ID>IN_0</ID>1611 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC2</lparam></gate>
<gate>
<ID>1498</ID>
<type>DE_TO</type>
<position>632.5,1391</position>
<input>
<ID>IN_0</ID>1566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>1499</ID>
<type>AE_SMALL_INVERTER</type>
<position>648.5,1388</position>
<input>
<ID>IN_0</ID>1567 </input>
<output>
<ID>OUT_0</ID>1568 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1500</ID>
<type>AE_SMALL_INVERTER</type>
<position>648.5,1382</position>
<input>
<ID>IN_0</ID>1568 </input>
<output>
<ID>OUT_0</ID>1569 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1501</ID>
<type>AE_SMALL_INVERTER</type>
<position>643,1380</position>
<input>
<ID>IN_0</ID>1569 </input>
<output>
<ID>OUT_0</ID>1570 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1502</ID>
<type>AE_SMALL_INVERTER</type>
<position>635,1380</position>
<input>
<ID>IN_0</ID>1570 </input>
<output>
<ID>OUT_0</ID>1572 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1503</ID>
<type>DE_TO</type>
<position>746.5,1489.5</position>
<input>
<ID>IN_0</ID>1612 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC3</lparam></gate>
<gate>
<ID>1504</ID>
<type>AE_OR2</type>
<position>633.5,1387</position>
<input>
<ID>IN_0</ID>1564 </input>
<input>
<ID>IN_1</ID>1572 </input>
<output>
<ID>OUT</ID>1571 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1505</ID>
<type>DE_TO</type>
<position>654.5,1390</position>
<input>
<ID>IN_0</ID>1567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1506</ID>
<type>FF_GND</type>
<position>741.5,1481.5</position>
<output>
<ID>OUT_0</ID>1615 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1507</ID>
<type>DE_TO</type>
<position>588.5,1506.5</position>
<input>
<ID>IN_0</ID>1573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Do step</lparam></gate>
<gate>
<ID>1508</ID>
<type>CC_PULSE</type>
<position>528.5,1389.5</position>
<output>
<ID>OUT_0</ID>1574 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1509</ID>
<type>DE_TO</type>
<position>538.5,1389.5</position>
<input>
<ID>IN_0</ID>1574 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Input</lparam></gate>
<gate>
<ID>1510</ID>
<type>DA_FROM</type>
<position>609,1392</position>
<input>
<ID>IN_0</ID>1618 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID rs</lparam></gate>
<gate>
<ID>1511</ID>
<type>DE_TO</type>
<position>737,1415</position>
<input>
<ID>IN_0</ID>1694 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACS</lparam></gate>
<gate>
<ID>1512</ID>
<type>DE_TO</type>
<position>737,1413</position>
<input>
<ID>IN_0</ID>1695 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MemClk</lparam></gate>
<gate>
<ID>1513</ID>
<type>DE_TO</type>
<position>737,1407</position>
<input>
<ID>IN_0</ID>1698 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCL</lparam></gate>
<gate>
<ID>1514</ID>
<type>DE_TO</type>
<position>737,1405</position>
<input>
<ID>IN_0</ID>1699 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDBR</lparam></gate>
<gate>
<ID>1515</ID>
<type>DE_TO</type>
<position>737,1411</position>
<input>
<ID>IN_0</ID>1696 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRS</lparam></gate>
<gate>
<ID>1516</ID>
<type>DE_TO</type>
<position>737,1409</position>
<input>
<ID>IN_0</ID>1697 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCS</lparam></gate>
<gate>
<ID>1517</ID>
<type>DE_TO</type>
<position>737,1399</position>
<input>
<ID>IN_0</ID>1702 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MemR</lparam></gate>
<gate>
<ID>1518</ID>
<type>DE_TO</type>
<position>737,1397</position>
<input>
<ID>IN_0</ID>1703 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MARW</lparam></gate>
<gate>
<ID>1519</ID>
<type>DE_TO</type>
<position>737,1391</position>
<input>
<ID>IN_0</ID>1706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACW1</lparam></gate>
<gate>
<ID>1520</ID>
<type>DE_TO</type>
<position>737,1389</position>
<input>
<ID>IN_0</ID>1707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond</lparam></gate>
<gate>
<ID>1521</ID>
<type>DE_TO</type>
<position>737,1395</position>
<input>
<ID>IN_0</ID>1704 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IRW</lparam></gate>
<gate>
<ID>1522</ID>
<type>DE_TO</type>
<position>737,1393</position>
<input>
<ID>IN_0</ID>1705 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW</lparam></gate>
<gate>
<ID>1523</ID>
<type>DE_TO</type>
<position>737,1403</position>
<input>
<ID>IN_0</ID>1700 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDBW</lparam></gate>
<gate>
<ID>1524</ID>
<type>BM_ROM_16x16</type>
<position>728,1436</position>
<input>
<ID>ADDRESS_0</ID>1708 </input>
<input>
<ID>ADDRESS_1</ID>1709 </input>
<input>
<ID>ADDRESS_10</ID>1740 </input>
<input>
<ID>ADDRESS_11</ID>1740 </input>
<input>
<ID>ADDRESS_12</ID>1740 </input>
<input>
<ID>ADDRESS_13</ID>1740 </input>
<input>
<ID>ADDRESS_14</ID>1740 </input>
<input>
<ID>ADDRESS_15</ID>1740 </input>
<input>
<ID>ADDRESS_2</ID>1710 </input>
<input>
<ID>ADDRESS_3</ID>1711 </input>
<input>
<ID>ADDRESS_4</ID>1712 </input>
<input>
<ID>ADDRESS_5</ID>1713 </input>
<input>
<ID>ADDRESS_6</ID>1714 </input>
<input>
<ID>ADDRESS_7</ID>1715 </input>
<input>
<ID>ADDRESS_8</ID>1740 </input>
<input>
<ID>ADDRESS_9</ID>1740 </input>
<output>
<ID>DATA_OUT_0</ID>1692 </output>
<output>
<ID>DATA_OUT_1</ID>1693 </output>
<output>
<ID>DATA_OUT_10</ID>1702 </output>
<output>
<ID>DATA_OUT_11</ID>1703 </output>
<output>
<ID>DATA_OUT_12</ID>1704 </output>
<output>
<ID>DATA_OUT_13</ID>1705 </output>
<output>
<ID>DATA_OUT_14</ID>1706 </output>
<output>
<ID>DATA_OUT_15</ID>1707 </output>
<output>
<ID>DATA_OUT_2</ID>1694 </output>
<output>
<ID>DATA_OUT_3</ID>1695 </output>
<output>
<ID>DATA_OUT_4</ID>1696 </output>
<output>
<ID>DATA_OUT_5</ID>1697 </output>
<output>
<ID>DATA_OUT_6</ID>1698 </output>
<output>
<ID>DATA_OUT_7</ID>1699 </output>
<output>
<ID>DATA_OUT_8</ID>1700 </output>
<output>
<ID>DATA_OUT_9</ID>1701 </output>
<input>
<ID>ENABLE_0</ID>1741 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 16</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 32</lparam>
<lparam>Address:1 2080</lparam>
<lparam>Address:2 1024</lparam>
<lparam>Address:3 5120</lparam>
<lparam>Address:4 32</lparam>
<lparam>Address:5 288</lparam>
<lparam>Address:6 16</lparam>
<lparam>Address:7 2064</lparam>
<lparam>Address:8 132</lparam>
<lparam>Address:9 140</lparam>
<lparam>Address:10 16</lparam>
<lparam>Address:11 16656</lparam>
<lparam>Address:12 16896</lparam>
<lparam>Address:13 130</lparam>
<lparam>Address:14 706</lparam>
<lparam>Address:15 8260</lparam>
<lparam>Address:16 32</lparam>
<lparam>Address:17 2080</lparam>
<lparam>Address:18 1024</lparam>
<lparam>Address:19 5120</lparam>
<lparam>Address:20 8192</lparam>
<lparam>Address:21 16</lparam>
<lparam>Address:22 2064</lparam>
<lparam>Address:23 1024</lparam>
<lparam>Address:24 1280</lparam>
<lparam>Address:25 512</lparam>
<lparam>Address:26 2</lparam>
<lparam>Address:27 1</lparam>
<lparam>Address:32 32</lparam>
<lparam>Address:33 2080</lparam>
<lparam>Address:34 1024</lparam>
<lparam>Address:35 5120</lparam>
<lparam>Address:36 8192</lparam>
<lparam>Address:37 16</lparam>
<lparam>Address:38 2064</lparam>
<lparam>Address:39 4</lparam>
<lparam>Address:40 12</lparam>
<lparam>Address:41 1</lparam>
<lparam>Address:48 32</lparam>
<lparam>Address:49 2080</lparam>
<lparam>Address:50 1024</lparam>
<lparam>Address:51 5120</lparam>
<lparam>Address:52 8192</lparam>
<lparam>Address:53 16</lparam>
<lparam>Address:54 2064</lparam>
<lparam>Address:55 1024</lparam>
<lparam>Address:56 1280</lparam>
<lparam>Address:57 512</lparam>
<lparam>Address:58 1</lparam>
<lparam>Address:64 32</lparam>
<lparam>Address:65 2080</lparam>
<lparam>Address:66 1024</lparam>
<lparam>Address:67 5120</lparam>
<lparam>Address:68 8192</lparam>
<lparam>Address:69 16</lparam>
<lparam>Address:70 2064</lparam>
<lparam>Address:71 1024</lparam>
<lparam>Address:72 1280</lparam>
<lparam>Address:73 512</lparam>
<lparam>Address:74 1</lparam>
<lparam>Address:80 32</lparam>
<lparam>Address:81 2080</lparam>
<lparam>Address:82 1024</lparam>
<lparam>Address:83 5120</lparam>
<lparam>Address:84 8192</lparam>
<lparam>Address:85 16</lparam>
<lparam>Address:86 2064</lparam>
<lparam>Address:87 1024</lparam>
<lparam>Address:88 1280</lparam>
<lparam>Address:89 384</lparam>
<lparam>Address:90 2176</lparam>
<lparam>Address:91 1280</lparam>
<lparam>Address:112 1</lparam>
<lparam>Address:128 32</lparam>
<lparam>Address:129 2080</lparam>
<lparam>Address:130 1024</lparam>
<lparam>Address:131 5120</lparam>
<lparam>Address:132 8192</lparam>
<lparam>Address:133 16</lparam>
<lparam>Address:134 2064</lparam>
<lparam>Address:135 32768</lparam>
<lparam>Address:136 1</lparam>
<lparam>Address:144 32</lparam>
<lparam>Address:145 2080</lparam>
<lparam>Address:146 1024</lparam>
<lparam>Address:147 5120</lparam>
<lparam>Address:148 80</lparam>
<lparam>Address:149 8272</lparam>
<lparam>Address:150 1</lparam>
<lparam>Address:160 32</lparam>
<lparam>Address:161 2080</lparam>
<lparam>Address:162 1024</lparam>
<lparam>Address:163 5120</lparam>
<lparam>Address:164 80</lparam>
<lparam>Address:165 2064</lparam>
<lparam>Address:166 4</lparam>
<lparam>Address:167 516</lparam>
<lparam>Address:168 1</lparam>
<lparam>Address:176 32</lparam>
<lparam>Address:177 2080</lparam>
<lparam>Address:178 1024</lparam>
<lparam>Address:179 5120</lparam>
<lparam>Address:180 8192</lparam>
<lparam>Address:181 2064</lparam>
<lparam>Address:182 1024</lparam>
<lparam>Address:183 1280</lparam>
<lparam>Address:184 384</lparam>
<lparam>Address:185 2176</lparam>
<lparam>Address:186 1024</lparam>
<lparam>Address:187 1280</lparam>
<lparam>Address:188 640</lparam>
<lparam>Address:189 1</lparam>
<lparam>Address:192 32</lparam>
<lparam>Address:193 2080</lparam>
<lparam>Address:194 1024</lparam>
<lparam>Address:195 5120</lparam>
<lparam>Address:196 8192</lparam>
<lparam>Address:197 16</lparam>
<lparam>Address:198 2064</lparam>
<lparam>Address:199 1024</lparam>
<lparam>Address:200 1280</lparam>
<lparam>Address:201 128</lparam>
<lparam>Address:202 8384</lparam>
<lparam>Address:203 1</lparam>
<lparam>Address:208 32</lparam>
<lparam>Address:209 2080</lparam>
<lparam>Address:210 1024</lparam>
<lparam>Address:211 5120</lparam>
<lparam>Address:212 8192</lparam>
<lparam>Address:213 16</lparam>
<lparam>Address:214 2064</lparam>
<lparam>Address:215 1280</lparam>
<lparam>Address:216 3072</lparam>
<lparam>Address:217 1280</lparam>
<lparam>Address:218 512</lparam>
<lparam>Address:219 1</lparam>
<lparam>Address:224 32</lparam>
<lparam>Address:225 2080</lparam>
<lparam>Address:226 1024</lparam>
<lparam>Address:227 5120</lparam>
<lparam>Address:228 8192</lparam>
<lparam>Address:229 16</lparam>
<lparam>Address:230 2064</lparam>
<lparam>Address:231 1280</lparam>
<lparam>Address:232 3072</lparam>
<lparam>Address:233 4</lparam>
<lparam>Address:234 12</lparam>
<lparam>Address:235 1</lparam></gate>
<gate>
<ID>1525</ID>
<type>DE_TO</type>
<position>737,1401</position>
<input>
<ID>IN_0</ID>1701 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACW</lparam></gate>
<gate>
<ID>1526</ID>
<type>AM_REGISTER16</type>
<position>599,1406.5</position>
<input>
<ID>IN_0</ID>1468 </input>
<input>
<ID>IN_1</ID>1461 </input>
<input>
<ID>IN_10</ID>1470 </input>
<input>
<ID>IN_11</ID>1458 </input>
<input>
<ID>IN_12</ID>1466 </input>
<input>
<ID>IN_13</ID>1459 </input>
<input>
<ID>IN_14</ID>1467 </input>
<input>
<ID>IN_15</ID>1460 </input>
<input>
<ID>IN_2</ID>1469 </input>
<input>
<ID>IN_3</ID>1462 </input>
<input>
<ID>IN_4</ID>1463 </input>
<input>
<ID>IN_5</ID>1416 </input>
<input>
<ID>IN_6</ID>1464 </input>
<input>
<ID>IN_7</ID>1456 </input>
<input>
<ID>IN_8</ID>1465 </input>
<input>
<ID>IN_9</ID>1457 </input>
<output>
<ID>OUT_0</ID>1602 </output>
<output>
<ID>OUT_1</ID>1594 </output>
<output>
<ID>OUT_10</ID>1597 </output>
<output>
<ID>OUT_11</ID>1590 </output>
<output>
<ID>OUT_12</ID>1596 </output>
<output>
<ID>OUT_13</ID>1589 </output>
<output>
<ID>OUT_14</ID>1595 </output>
<output>
<ID>OUT_15</ID>1588 </output>
<output>
<ID>OUT_2</ID>1601 </output>
<output>
<ID>OUT_3</ID>1593 </output>
<output>
<ID>OUT_4</ID>1600 </output>
<output>
<ID>OUT_5</ID>1592 </output>
<output>
<ID>OUT_6</ID>1599 </output>
<output>
<ID>OUT_7</ID>1591 </output>
<output>
<ID>OUT_8</ID>1598 </output>
<output>
<ID>OUT_9</ID>1587 </output>
<output>
<ID>carry_out</ID>1490 </output>
<input>
<ID>clear</ID>1618 </input>
<input>
<ID>clock</ID>1614 </input>
<input>
<ID>count_enable</ID>1487 </input>
<input>
<ID>count_up</ID>1489 </input>
<input>
<ID>load</ID>1488 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1527</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>608.5,1406.5</position>
<input>
<ID>ENABLE_0</ID>1603 </input>
<input>
<ID>IN_0</ID>1602 </input>
<input>
<ID>IN_1</ID>1594 </input>
<input>
<ID>IN_10</ID>1597 </input>
<input>
<ID>IN_11</ID>1590 </input>
<input>
<ID>IN_12</ID>1596 </input>
<input>
<ID>IN_13</ID>1589 </input>
<input>
<ID>IN_14</ID>1595 </input>
<input>
<ID>IN_15</ID>1588 </input>
<input>
<ID>IN_2</ID>1601 </input>
<input>
<ID>IN_3</ID>1593 </input>
<input>
<ID>IN_4</ID>1600 </input>
<input>
<ID>IN_5</ID>1592 </input>
<input>
<ID>IN_6</ID>1599 </input>
<input>
<ID>IN_7</ID>1591 </input>
<input>
<ID>IN_8</ID>1598 </input>
<input>
<ID>IN_9</ID>1587 </input>
<output>
<ID>OUT_0</ID>1473 </output>
<output>
<ID>OUT_1</ID>1486 </output>
<output>
<ID>OUT_10</ID>1478 </output>
<output>
<ID>OUT_11</ID>1481 </output>
<output>
<ID>OUT_12</ID>1471 </output>
<output>
<ID>OUT_13</ID>1482 </output>
<output>
<ID>OUT_14</ID>1472 </output>
<output>
<ID>OUT_15</ID>1483 </output>
<output>
<ID>OUT_2</ID>1474 </output>
<output>
<ID>OUT_3</ID>1485 </output>
<output>
<ID>OUT_4</ID>1475 </output>
<output>
<ID>OUT_5</ID>1484 </output>
<output>
<ID>OUT_6</ID>1476 </output>
<output>
<ID>OUT_7</ID>1479 </output>
<output>
<ID>OUT_8</ID>1477 </output>
<output>
<ID>OUT_9</ID>1480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1528</ID>
<type>DA_FROM</type>
<position>608.5,1421</position>
<input>
<ID>IN_0</ID>1603 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID PCS</lparam></gate>
<gate>
<ID>1529</ID>
<type>DA_FROM</type>
<position>710.5,1420.5</position>
<input>
<ID>IN_0</ID>1708 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>1530</ID>
<type>DA_FROM</type>
<position>710.5,1423</position>
<input>
<ID>IN_0</ID>1709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>1531</ID>
<type>DA_FROM</type>
<position>710.5,1425.5</position>
<input>
<ID>IN_0</ID>1710 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>1532</ID>
<type>DA_FROM</type>
<position>710.5,1428</position>
<input>
<ID>IN_0</ID>1711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>1533</ID>
<type>DA_FROM</type>
<position>710.5,1430.5</position>
<input>
<ID>IN_0</ID>1712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC0</lparam></gate>
<gate>
<ID>1534</ID>
<type>DA_FROM</type>
<position>710,1435</position>
<input>
<ID>IN_0</ID>1714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC2</lparam></gate>
<gate>
<ID>1535</ID>
<type>DA_FROM</type>
<position>710.5,1432.5</position>
<input>
<ID>IN_0</ID>1713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC1</lparam></gate>
<gate>
<ID>1536</ID>
<type>DA_FROM</type>
<position>710,1437.5</position>
<input>
<ID>IN_0</ID>1715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OC3</lparam></gate>
<gate>
<ID>1537</ID>
<type>AA_REGISTER4</type>
<position>751.5,1436.5</position>
<output>
<ID>OUT_0</ID>1719 </output>
<output>
<ID>OUT_1</ID>1718 </output>
<output>
<ID>OUT_2</ID>1717 </output>
<output>
<ID>OUT_3</ID>1716 </output>
<input>
<ID>clear</ID>1725 </input>
<input>
<ID>clock</ID>1724 </input>
<input>
<ID>count_enable</ID>1720 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1538</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1471.5,685,1471.5</points>
<connection>
<GID>1453</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_8</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1471.5,673,1490</points>
<intersection>1471.5 0</intersection>
<intersection>1490 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1490,684,1490</points>
<connection>
<GID>1281</GID>
<name>IN_8</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>1539</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1469.5,685,1469.5</points>
<connection>
<GID>1454</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_6</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1469.5,673,1488</points>
<intersection>1469.5 0</intersection>
<intersection>1488 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1488,684,1488</points>
<connection>
<GID>1281</GID>
<name>IN_6</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>1540</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1467.5,685,1467.5</points>
<connection>
<GID>1455</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_4</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1467.5,673,1486</points>
<intersection>1467.5 0</intersection>
<intersection>1486 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1486,684,1486</points>
<connection>
<GID>1281</GID>
<name>IN_4</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>1541</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1465.5,685,1465.5</points>
<connection>
<GID>1456</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_2</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1465.5,673,1484</points>
<intersection>1465.5 0</intersection>
<intersection>1484 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1484,684,1484</points>
<connection>
<GID>1281</GID>
<name>IN_2</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>513.5,1517,513.5,1521</points>
<connection>
<GID>2</GID>
<name>count_up</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1542</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1463.5,685,1463.5</points>
<connection>
<GID>1457</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_0</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1463.5,673,1482</points>
<intersection>1463.5 0</intersection>
<intersection>1482 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1482,684,1482</points>
<connection>
<GID>1281</GID>
<name>IN_0</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514.5,1488,514.5,1498</points>
<intersection>1488 1</intersection>
<intersection>1498 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>508,1488,514.5,1488</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>510.5 4</intersection>
<intersection>514.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>513.5,1498,514.5,1498</points>
<connection>
<GID>2</GID>
<name>clear</name></connection>
<intersection>514.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>510.5,1488,510.5,1491</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>1488 1</intersection></vsegment></shape></wire>
<wire>
<ID>1543</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1477.5,748,1477.5</points>
<connection>
<GID>1464</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1426</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>511.5,1497,511.5,1498</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>1544</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1463.5,748,1463.5</points>
<connection>
<GID>1464</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1461</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,1489.5,512.5,1491</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>1489.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512.5,1489.5,526,1489.5</points>
<intersection>512.5 0</intersection>
<intersection>526 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>526,1489.5,526,1505.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>1489.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1545</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1465.5,748,1465.5</points>
<connection>
<GID>1464</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>731,1501,734.5,1501</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1546</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1467.5,748,1467.5</points>
<connection>
<GID>1464</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1459</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>512.5,1517,512.5,1520.5</points>
<connection>
<GID>2</GID>
<name>count_enable</name></connection>
<intersection>1520.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>512.5,1520.5,516.5,1520.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>512.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1547</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1469.5,748,1469.5</points>
<connection>
<GID>1464</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1430</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>522.5,1521.5,524,1521.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1548</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1471.5,748,1471.5</points>
<connection>
<GID>1464</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1429</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,1511.5,579,1520.5</points>
<intersection>1511.5 1</intersection>
<intersection>1520.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>579,1511.5,725,1511.5</points>
<intersection>579 0</intersection>
<intersection>725 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>522.5,1520.5,579,1520.5</points>
<intersection>522.5 7</intersection>
<intersection>579 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>725,1504,725,1511.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>1511.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>522.5,1519.5,522.5,1520.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>1520.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>1549</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1473.5,748,1473.5</points>
<connection>
<GID>1464</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1428</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1550</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1470.5,755.5,1470.5</points>
<connection>
<GID>1464</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1422</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1551</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1472.5,755.5,1472.5</points>
<connection>
<GID>1464</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1552</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1474.5,755.5,1474.5</points>
<connection>
<GID>1464</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1420</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1553</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1476.5,755.5,1476.5</points>
<connection>
<GID>1464</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1419</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1554</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1478.5,755.5,1478.5</points>
<connection>
<GID>1464</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1418</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1555</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1468.5,755.5,1468.5</points>
<connection>
<GID>1464</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1466.5,755.5,1466.5</points>
<connection>
<GID>1464</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1424</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1557</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1464.5,755.5,1464.5</points>
<connection>
<GID>1464</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1425</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667,1457.5,667,1461.5</points>
<connection>
<GID>1458</GID>
<name>clock</name></connection>
<intersection>1457.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>665.5,1457.5,667,1457.5</points>
<connection>
<GID>1468</GID>
<name>OUT</name></connection>
<intersection>667 0</intersection></hsegment></shape></wire>
<wire>
<ID>1559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>656.5,1458.5,659.5,1458.5</points>
<connection>
<GID>1473</GID>
<name>IN_0</name></connection>
<connection>
<GID>1468</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1560</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>656.5,1456.5,659.5,1456.5</points>
<connection>
<GID>1477</GID>
<name>IN_0</name></connection>
<connection>
<GID>1468</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1561</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>669,1457.5,669,1461.5</points>
<connection>
<GID>1458</GID>
<name>clear</name></connection>
<intersection>1457.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>669,1457.5,670.5,1457.5</points>
<connection>
<GID>1436</GID>
<name>IN_0</name></connection>
<intersection>669 0</intersection></hsegment></shape></wire>
<wire>
<ID>1562</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>530.5,1407,536.5,1407</points>
<connection>
<GID>1482</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1489</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1563</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>636.5,1393,645.5,1393</points>
<intersection>636.5 5</intersection>
<intersection>645.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>645.5,1387,645.5,1393</points>
<intersection>1387 8</intersection>
<intersection>1393 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>636.5,1390,636.5,1393</points>
<intersection>1390 9</intersection>
<intersection>1393 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>644,1387,645.5,1387</points>
<connection>
<GID>1491</GID>
<name>OUTINV_0</name></connection>
<intersection>645.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>636.5,1390,638,1390</points>
<connection>
<GID>1491</GID>
<name>IN_0</name></connection>
<intersection>636.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>619,1388,630.5,1388</points>
<connection>
<GID>1493</GID>
<name>IN_0</name></connection>
<connection>
<GID>1504</GID>
<name>IN_0</name></connection>
<intersection>620.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>620.5,1388,620.5,1391</points>
<intersection>1388 1</intersection>
<intersection>1391 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>620.5,1391,621.5,1391</points>
<connection>
<GID>1495</GID>
<name>IN_0</name></connection>
<intersection>620.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>1565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>625.5,1391,626.5,1391</points>
<connection>
<GID>1495</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1496</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>630.5,1391,630.5,1391</points>
<connection>
<GID>1496</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1498</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1567</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>644,1390,652.5,1390</points>
<connection>
<GID>1499</GID>
<name>IN_0</name></connection>
<connection>
<GID>1491</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1505</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>648.5,1384,648.5,1386</points>
<connection>
<GID>1500</GID>
<name>IN_0</name></connection>
<connection>
<GID>1499</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1569</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>645,1380,648.5,1380</points>
<connection>
<GID>1500</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1501</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1570</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>637,1380,641,1380</points>
<connection>
<GID>1502</GID>
<name>IN_0</name></connection>
<connection>
<GID>1501</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1571</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>636.5,1387,638,1387</points>
<connection>
<GID>1504</GID>
<name>OUT</name></connection>
<connection>
<GID>1491</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1572</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>629,1380,629,1386</points>
<intersection>1380 2</intersection>
<intersection>1386 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>629,1386,630.5,1386</points>
<connection>
<GID>1504</GID>
<name>IN_1</name></connection>
<intersection>629 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>629,1380,633,1380</points>
<connection>
<GID>1502</GID>
<name>OUT_0</name></connection>
<intersection>629 0</intersection></hsegment></shape></wire>
<wire>
<ID>1573</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>584.5,1506.5,586.5,1506.5</points>
<connection>
<GID>1208</GID>
<name>OUT</name></connection>
<connection>
<GID>1507</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1574</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>530.5,1389.5,536.5,1389.5</points>
<connection>
<GID>1508</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1509</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1575</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1472.5,741.5,1472.5</points>
<connection>
<GID>1463</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1464</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1576</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1474.5,741.5,1474.5</points>
<connection>
<GID>1463</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1464</GID>
<name>IN_11</name></connection>
<intersection>740 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>740,1474.5,740,1496.5</points>
<intersection>1474.5 1</intersection>
<intersection>1496.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>740,1496.5,745,1496.5</points>
<connection>
<GID>1211</GID>
<name>IN_0</name></connection>
<intersection>740 2</intersection></hsegment></shape></wire>
<wire>
<ID>1577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1470.5,741.5,1470.5</points>
<connection>
<GID>1463</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1464</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1578</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1468.5,741.5,1468.5</points>
<connection>
<GID>1463</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1464</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1579</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1466.5,741.5,1466.5</points>
<connection>
<GID>1463</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1464</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>736,1464.5,741.5,1464.5</points>
<connection>
<GID>1463</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1464</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1581</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1473.5,741.5,1473.5</points>
<connection>
<GID>1463</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1464</GID>
<name>IN_10</name></connection>
<intersection>740.5 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>740.5,1473.5,740.5,1494</points>
<intersection>1473.5 0</intersection>
<intersection>1494 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>740.5,1494,745,1494</points>
<connection>
<GID>1212</GID>
<name>IN_0</name></connection>
<intersection>740.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>1582</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1471.5,741.5,1471.5</points>
<connection>
<GID>1463</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1464</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1583</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1469.5,741.5,1469.5</points>
<connection>
<GID>1463</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1464</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1584</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1467.5,741.5,1467.5</points>
<connection>
<GID>1463</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1464</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1585</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1465.5,741.5,1465.5</points>
<connection>
<GID>1463</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1464</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1586</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>736,1463.5,741.5,1463.5</points>
<connection>
<GID>1463</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1464</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1587</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1408,606.5,1408</points>
<connection>
<GID>1526</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1527</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1588</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1414,606.5,1414</points>
<connection>
<GID>1526</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1527</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1589</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1412,606.5,1412</points>
<connection>
<GID>1526</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1527</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1410,606.5,1410</points>
<connection>
<GID>1526</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1527</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1591</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1406,606.5,1406</points>
<connection>
<GID>1526</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1527</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1592</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1404,606.5,1404</points>
<connection>
<GID>1526</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1527</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1593</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1402,606.5,1402</points>
<connection>
<GID>1526</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1527</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1594</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>604,1400,606.5,1400</points>
<connection>
<GID>1526</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1527</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1595</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1413,606.5,1413</points>
<connection>
<GID>1526</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1527</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1596</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1411,606.5,1411</points>
<connection>
<GID>1526</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1527</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1597</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1409,606.5,1409</points>
<connection>
<GID>1526</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1527</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1598</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1407,606.5,1407</points>
<connection>
<GID>1526</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1527</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1599</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1405,606.5,1405</points>
<connection>
<GID>1526</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1527</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1600</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1403,606.5,1403</points>
<connection>
<GID>1526</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1527</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1601</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1401,606.5,1401</points>
<connection>
<GID>1526</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1527</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1602</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>604,1399,606.5,1399</points>
<connection>
<GID>1526</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1527</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1603</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>608.5,1415.5,608.5,1419</points>
<connection>
<GID>1527</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1528</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>729,1456.5,730,1456.5</points>
<connection>
<GID>1466</GID>
<name>OUT</name></connection>
<intersection>730 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>730,1456.5,730,1461.5</points>
<connection>
<GID>1463</GID>
<name>clock</name></connection>
<intersection>1456.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1605</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>722,1455.5,723,1455.5</points>
<connection>
<GID>1467</GID>
<name>IN_0</name></connection>
<connection>
<GID>1466</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1606</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>732,1456.5,732,1461.5</points>
<connection>
<GID>1462</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>1607</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>743.5,1480,743.5,1481.5</points>
<connection>
<GID>1464</GID>
<name>ENABLE_0</name></connection>
<intersection>1481.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>743.5,1481.5,747,1481.5</points>
<connection>
<GID>1465</GID>
<name>IN_0</name></connection>
<intersection>743.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1608</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>730,1480.5,730,1482.5</points>
<connection>
<GID>1463</GID>
<name>load</name></connection>
<connection>
<GID>1488</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1609</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>738.5,1475.5,738.5,1507</points>
<intersection>1475.5 1</intersection>
<intersection>1483.5 2</intersection>
<intersection>1507 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>736,1475.5,738.5,1475.5</points>
<connection>
<GID>1463</GID>
<name>OUT_12</name></connection>
<intersection>738.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>738.5,1483.5,744.5,1483.5</points>
<connection>
<GID>1492</GID>
<name>IN_0</name></connection>
<intersection>738.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>731,1507,738.5,1507</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>738.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>738,1476.5,738,1505</points>
<intersection>1476.5 1</intersection>
<intersection>1485.5 2</intersection>
<intersection>1505 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>736,1476.5,738,1476.5</points>
<connection>
<GID>1463</GID>
<name>OUT_13</name></connection>
<intersection>738 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>738,1485.5,744.5,1485.5</points>
<connection>
<GID>1494</GID>
<name>IN_0</name></connection>
<intersection>738 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>731,1505,738,1505</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>738 0</intersection></hsegment></shape></wire>
<wire>
<ID>1611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>737.5,1477.5,737.5,1503</points>
<intersection>1477.5 1</intersection>
<intersection>1487.5 2</intersection>
<intersection>1503 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>736,1477.5,737.5,1477.5</points>
<connection>
<GID>1463</GID>
<name>OUT_14</name></connection>
<intersection>737.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>737.5,1487.5,744.5,1487.5</points>
<connection>
<GID>1497</GID>
<name>IN_0</name></connection>
<intersection>737.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>731,1503,737.5,1503</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>737.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>737,1478.5,737,1497</points>
<intersection>1478.5 1</intersection>
<intersection>1489.5 2</intersection>
<intersection>1497 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>736,1478.5,737,1478.5</points>
<connection>
<GID>1463</GID>
<name>OUT_15</name></connection>
<intersection>737 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>737,1489.5,744.5,1489.5</points>
<connection>
<GID>1503</GID>
<name>IN_0</name></connection>
<intersection>737 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>734.5,1497,737,1497</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>737 0</intersection></hsegment></shape></wire>
<wire>
<ID>1613</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>720,1457.5,723,1457.5</points>
<connection>
<GID>1470</GID>
<name>IN_0</name></connection>
<connection>
<GID>1466</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1614</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>598,1390,598,1397</points>
<connection>
<GID>1545</GID>
<name>OUT</name></connection>
<connection>
<GID>1526</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>1615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>741.5,1475.5,741.5,1480.5</points>
<connection>
<GID>1464</GID>
<name>IN_15</name></connection>
<connection>
<GID>1464</GID>
<name>IN_14</name></connection>
<connection>
<GID>1464</GID>
<name>IN_13</name></connection>
<connection>
<GID>1464</GID>
<name>IN_12</name></connection>
<connection>
<GID>1506</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1616</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>678,1430,685.5,1430</points>
<connection>
<GID>1562</GID>
<name>write_clock</name></connection>
<connection>
<GID>1260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1617</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>587.5,1384,592,1384</points>
<connection>
<GID>1554</GID>
<name>IN_0</name></connection>
<intersection>592 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>592,1384,592,1389</points>
<connection>
<GID>1545</GID>
<name>IN_1</name></connection>
<intersection>1384 0</intersection></vsegment></shape></wire>
<wire>
<ID>1618</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600,1392,600,1397</points>
<connection>
<GID>1526</GID>
<name>clear</name></connection>
<intersection>1392 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>600,1392,607,1392</points>
<connection>
<GID>1510</GID>
<name>IN_0</name></connection>
<intersection>600 0</intersection></hsegment></shape></wire>
<wire>
<ID>1619</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>588.5,1391,592,1391</points>
<connection>
<GID>1557</GID>
<name>OUT</name></connection>
<connection>
<GID>1545</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1620</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>581.5,1394,581.5,1394</points>
<connection>
<GID>1550</GID>
<name>IN_0</name></connection>
<connection>
<GID>1557</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1621</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>581.5,1392,581.5,1392</points>
<connection>
<GID>1557</GID>
<name>IN_1</name></connection>
<connection>
<GID>1558</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1622</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>581.5,1390,581.5,1390</points>
<connection>
<GID>1557</GID>
<name>IN_2</name></connection>
<connection>
<GID>1559</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1623</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>580,1388,581.5,1388</points>
<connection>
<GID>1560</GID>
<name>IN_0</name></connection>
<connection>
<GID>1557</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1624</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1421,660,1421</points>
<connection>
<GID>1564</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1422,660,1422</points>
<connection>
<GID>1564</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1626</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1423,660,1423</points>
<connection>
<GID>1564</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1627</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1424,660,1424</points>
<connection>
<GID>1564</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1628</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1425,660,1425</points>
<connection>
<GID>1564</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1629</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1426,660,1426</points>
<connection>
<GID>1564</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1630</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1427,660,1427</points>
<connection>
<GID>1564</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1631</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1428,660,1428</points>
<connection>
<GID>1564</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1632</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1429,660,1429</points>
<connection>
<GID>1564</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1633</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1430,660,1430</points>
<connection>
<GID>1564</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1634</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1431,660,1431</points>
<connection>
<GID>1564</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1635</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1432,660,1432</points>
<connection>
<GID>1564</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1433,660,1433</points>
<connection>
<GID>1564</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1637</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1434,660,1434</points>
<connection>
<GID>1564</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1638</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1435,660,1435</points>
<connection>
<GID>1564</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1639</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1436,660,1436</points>
<connection>
<GID>1564</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1562</GID>
<name>ADDRESS_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>649.5,1416.5,649.5,1419</points>
<connection>
<GID>1564</GID>
<name>clock</name></connection>
<intersection>1416.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>649,1416.5,649.5,1416.5</points>
<connection>
<GID>1566</GID>
<name>OUT</name></connection>
<intersection>649.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1641</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>640,1417.5,643,1417.5</points>
<connection>
<GID>1568</GID>
<name>IN_0</name></connection>
<connection>
<GID>1566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1642</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>643,1415.5,643,1415.5</points>
<connection>
<GID>1566</GID>
<name>IN_1</name></connection>
<connection>
<GID>1569</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1643</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>676.5,1408.5,676.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_0</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1417 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>676.5,1417,703,1417</points>
<intersection>676.5 0</intersection>
<intersection>703 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>703,1408,703,1417</points>
<connection>
<GID>1572</GID>
<name>OUT_0</name></connection>
<intersection>1417 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>676,1408.5,676.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_15</name></connection>
<intersection>676.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1644</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>675.5,1408.5,675.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_1</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1416.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>675.5,1416.5,702,1416.5</points>
<intersection>675.5 0</intersection>
<intersection>702 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>702,1408,702,1416.5</points>
<connection>
<GID>1572</GID>
<name>OUT_1</name></connection>
<intersection>1416.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>675,1408.5,675.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_14</name></connection>
<intersection>675.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1645</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>674.5,1408.5,674.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_2</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1416 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>674.5,1416,701,1416</points>
<intersection>674.5 0</intersection>
<intersection>701 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>701,1408,701,1416</points>
<connection>
<GID>1572</GID>
<name>OUT_2</name></connection>
<intersection>1416 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>674,1408.5,674.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_13</name></connection>
<intersection>674.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1646</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673.5,1408.5,673.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_3</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1415.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>673.5,1415.5,700,1415.5</points>
<intersection>673.5 0</intersection>
<intersection>700 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>700,1408,700,1415.5</points>
<connection>
<GID>1572</GID>
<name>OUT_3</name></connection>
<intersection>1415.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>673,1408.5,673.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_12</name></connection>
<intersection>673.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672.5,1408.5,672.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_4</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1415 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>672.5,1415,699,1415</points>
<intersection>672.5 0</intersection>
<intersection>699 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>699,1408,699,1415</points>
<connection>
<GID>1572</GID>
<name>OUT_4</name></connection>
<intersection>1415 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>672,1408.5,672.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_11</name></connection>
<intersection>672.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>671.5,1408.5,671.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_5</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1414.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>671.5,1414.5,698,1414.5</points>
<intersection>671.5 0</intersection>
<intersection>698 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>698,1408,698,1414.5</points>
<connection>
<GID>1572</GID>
<name>OUT_5</name></connection>
<intersection>1414.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>671,1408.5,671.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_10</name></connection>
<intersection>671.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>670.5,1408.5,670.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_6</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1414 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>670.5,1414,697,1414</points>
<intersection>670.5 0</intersection>
<intersection>697 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>697,1408,697,1414</points>
<connection>
<GID>1572</GID>
<name>OUT_6</name></connection>
<intersection>1414 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>670,1408.5,670.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_9</name></connection>
<intersection>670.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1650</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>669.5,1408.5,669.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_7</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1413.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>669.5,1413.5,696,1413.5</points>
<intersection>669.5 0</intersection>
<intersection>696 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>696,1408,696,1413.5</points>
<connection>
<GID>1572</GID>
<name>OUT_7</name></connection>
<intersection>1413.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>669,1408.5,669.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_8</name></connection>
<intersection>669.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1651</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668.5,1408.5,668.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_8</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1413 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>668.5,1413,695,1413</points>
<intersection>668.5 0</intersection>
<intersection>695 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>695,1408,695,1413</points>
<connection>
<GID>1572</GID>
<name>OUT_8</name></connection>
<intersection>1413 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>668,1408.5,668.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_7</name></connection>
<intersection>668.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1652</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667.5,1408.5,667.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_9</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1412.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>667.5,1412.5,694,1412.5</points>
<intersection>667.5 0</intersection>
<intersection>694 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>694,1408,694,1412.5</points>
<connection>
<GID>1572</GID>
<name>OUT_9</name></connection>
<intersection>1412.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>667,1408.5,667.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_6</name></connection>
<intersection>667.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1653</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666.5,1408.5,666.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_10</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1412 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>666.5,1412,693,1412</points>
<intersection>666.5 0</intersection>
<intersection>693 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>693,1408,693,1412</points>
<connection>
<GID>1572</GID>
<name>OUT_10</name></connection>
<intersection>1412 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>666,1408.5,666.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_5</name></connection>
<intersection>666.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1654</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665.5,1408.5,665.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_11</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1411.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>665.5,1411.5,692,1411.5</points>
<intersection>665.5 0</intersection>
<intersection>692 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>692,1408,692,1411.5</points>
<connection>
<GID>1572</GID>
<name>OUT_11</name></connection>
<intersection>1411.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>665,1408.5,665.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_4</name></connection>
<intersection>665.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,1408.5,664.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_12</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1411 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>664.5,1411,691,1411</points>
<intersection>664.5 0</intersection>
<intersection>691 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>691,1408,691,1411</points>
<connection>
<GID>1572</GID>
<name>OUT_12</name></connection>
<intersection>1411 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>664,1408.5,664.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_3</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1656</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>663.5,1408.5,663.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_13</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1410.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>663.5,1410.5,690,1410.5</points>
<intersection>663.5 0</intersection>
<intersection>690 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>690,1408,690,1410.5</points>
<connection>
<GID>1572</GID>
<name>OUT_13</name></connection>
<intersection>1410.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>663,1408.5,663.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_2</name></connection>
<intersection>663.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1657</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>662.5,1408.5,662.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_14</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1410 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>662.5,1410,689,1410</points>
<intersection>662.5 0</intersection>
<intersection>689 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>689,1408,689,1410</points>
<connection>
<GID>1572</GID>
<name>OUT_14</name></connection>
<intersection>1410 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>662,1408.5,662.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_1</name></connection>
<intersection>662.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1658</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>661.5,1408.5,661.5,1417.5</points>
<connection>
<GID>1562</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>1562</GID>
<name>DATA_IN_15</name></connection>
<intersection>1408.5 21</intersection>
<intersection>1409.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>661.5,1409.5,688,1409.5</points>
<intersection>661.5 0</intersection>
<intersection>688 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>688,1408,688,1409.5</points>
<connection>
<GID>1572</GID>
<name>OUT_15</name></connection>
<intersection>1409.5 18</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>661,1408.5,661.5,1408.5</points>
<connection>
<GID>1571</GID>
<name>IN_0</name></connection>
<intersection>661.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1659</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>675,1396.5,675,1404.5</points>
<connection>
<GID>1580</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_14</name></connection></vsegment></shape></wire>
<wire>
<ID>1660</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>673,1396.5,673,1404.5</points>
<connection>
<GID>1579</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_12</name></connection></vsegment></shape></wire>
<wire>
<ID>1661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>671,1396.5,671,1404.5</points>
<connection>
<GID>1578</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_10</name></connection></vsegment></shape></wire>
<wire>
<ID>1662</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>669,1396.5,669,1404.5</points>
<connection>
<GID>1577</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_8</name></connection></vsegment></shape></wire>
<wire>
<ID>1663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667,1396.5,667,1404.5</points>
<connection>
<GID>1576</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_6</name></connection></vsegment></shape></wire>
<wire>
<ID>1664</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>665,1396.5,665,1404.5</points>
<connection>
<GID>1575</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_4</name></connection></vsegment></shape></wire>
<wire>
<ID>1665</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>663,1396.5,663,1404.5</points>
<connection>
<GID>1574</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>661,1396.5,661,1404.5</points>
<connection>
<GID>1573</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1667</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>688,1394,688,1404</points>
<connection>
<GID>1581</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>1668</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>692,1394,692,1404</points>
<connection>
<GID>1583</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>1669</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,1394,690,1404</points>
<connection>
<GID>1582</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>1670</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>694,1394,694,1404</points>
<connection>
<GID>1584</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>1671</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>696,1394,696,1404</points>
<connection>
<GID>1585</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>1672</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,1394,698,1404</points>
<connection>
<GID>1586</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>1673</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>700,1394,700,1404</points>
<connection>
<GID>1587</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>1674</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>702,1394,702,1404</points>
<connection>
<GID>1588</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1675</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>703,1401.5,703,1404</points>
<connection>
<GID>1596</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1676</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>701,1401.5,701,1404</points>
<connection>
<GID>1595</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>1677</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>699,1401.5,699,1404</points>
<connection>
<GID>1594</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>1678</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>697,1401.5,697,1404</points>
<connection>
<GID>1593</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>1679</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>695,1401.5,695,1404</points>
<connection>
<GID>1592</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>1680</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>693,1401.5,693,1404</points>
<connection>
<GID>1591</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>1681</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>691,1401.5,691,1404</points>
<connection>
<GID>1590</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>1682</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>689,1401.5,689,1404</points>
<connection>
<GID>1589</GID>
<name>IN_0</name></connection>
<connection>
<GID>1572</GID>
<name>IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>1683</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>662,1403.5,662,1404.5</points>
<connection>
<GID>1597</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>1684</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664,1403.5,664,1404.5</points>
<connection>
<GID>1598</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>1685</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>666,1403.5,666,1404.5</points>
<connection>
<GID>1599</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>1686</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>668,1403.5,668,1404.5</points>
<connection>
<GID>1600</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>1687</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>670,1403.5,670,1404.5</points>
<connection>
<GID>1601</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_9</name></connection></vsegment></shape></wire>
<wire>
<ID>1688</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>672,1403.5,672,1404.5</points>
<connection>
<GID>1602</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_11</name></connection></vsegment></shape></wire>
<wire>
<ID>1689</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>674,1403.5,674,1404.5</points>
<connection>
<GID>1603</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_13</name></connection></vsegment></shape></wire>
<wire>
<ID>1690</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>676,1403.5,676,1404.5</points>
<connection>
<GID>1604</GID>
<name>IN_0</name></connection>
<connection>
<GID>1571</GID>
<name>OUT_15</name></connection></vsegment></shape></wire>
<wire>
<ID>1691</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>651.5,1415.5,651.5,1419</points>
<connection>
<GID>1564</GID>
<name>clear</name></connection>
<intersection>1415.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>651.5,1415.5,652.5,1415.5</points>
<connection>
<GID>1606</GID>
<name>IN_0</name></connection>
<intersection>651.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1692</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>735.5,1419,735.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_0</name></connection>
<intersection>1419 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>735,1419,735.5,1419</points>
<connection>
<GID>1617</GID>
<name>IN_0</name></connection>
<intersection>735.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1693</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>734.5,1417,734.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_1</name></connection>
<intersection>1417 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>734.5,1417,735,1417</points>
<connection>
<GID>1618</GID>
<name>IN_0</name></connection>
<intersection>734.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>733.5,1415,733.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_2</name></connection>
<intersection>1415 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>733.5,1415,735,1415</points>
<connection>
<GID>1511</GID>
<name>IN_0</name></connection>
<intersection>733.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1695</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>732.5,1413,732.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_3</name></connection>
<intersection>1413 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>732.5,1413,735,1413</points>
<connection>
<GID>1512</GID>
<name>IN_0</name></connection>
<intersection>732.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>731.5,1411,731.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_4</name></connection>
<intersection>1411 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>731.5,1411,735,1411</points>
<connection>
<GID>1515</GID>
<name>IN_0</name></connection>
<intersection>731.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1697</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>730.5,1409,730.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_5</name></connection>
<intersection>1409 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>730.5,1409,735,1409</points>
<connection>
<GID>1516</GID>
<name>IN_0</name></connection>
<intersection>730.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1698</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>729.5,1407,729.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_6</name></connection>
<intersection>1407 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>729.5,1407,735,1407</points>
<connection>
<GID>1513</GID>
<name>IN_0</name></connection>
<intersection>729.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>728.5,1405,728.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_7</name></connection>
<intersection>1405 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>728.5,1405,735,1405</points>
<connection>
<GID>1514</GID>
<name>IN_0</name></connection>
<intersection>728.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1700</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>727.5,1403,727.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_8</name></connection>
<intersection>1403 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>727.5,1403,735,1403</points>
<connection>
<GID>1523</GID>
<name>IN_0</name></connection>
<intersection>727.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>726.5,1401,726.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_9</name></connection>
<intersection>1401 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>726.5,1401,735,1401</points>
<connection>
<GID>1525</GID>
<name>IN_0</name></connection>
<intersection>726.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1702</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>725.5,1399,725.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_10</name></connection>
<intersection>1399 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>725.5,1399,735,1399</points>
<connection>
<GID>1517</GID>
<name>IN_0</name></connection>
<intersection>725.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1703</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>724.5,1397,724.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_11</name></connection>
<intersection>1397 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>724.5,1397,735,1397</points>
<connection>
<GID>1518</GID>
<name>IN_0</name></connection>
<intersection>724.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>723.5,1395,723.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_12</name></connection>
<intersection>1395 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>723.5,1395,735,1395</points>
<connection>
<GID>1521</GID>
<name>IN_0</name></connection>
<intersection>723.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>722.5,1393,722.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_13</name></connection>
<intersection>1393 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>722.5,1393,735,1393</points>
<connection>
<GID>1522</GID>
<name>IN_0</name></connection>
<intersection>722.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1706</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>721.5,1391,721.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_14</name></connection>
<intersection>1391 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>721.5,1391,735,1391</points>
<connection>
<GID>1519</GID>
<name>IN_0</name></connection>
<intersection>721.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1707</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>720.5,1389,720.5,1425</points>
<connection>
<GID>1524</GID>
<name>DATA_OUT_15</name></connection>
<intersection>1389 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>720.5,1389,735,1389</points>
<connection>
<GID>1520</GID>
<name>IN_0</name></connection>
<intersection>720.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1708</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>718.5,1428.5,719,1428.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_0</name></connection>
<intersection>718.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>718.5,1420.5,718.5,1428.5</points>
<intersection>1420.5 21</intersection>
<intersection>1428.5 15</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712.5,1420.5,718.5,1420.5</points>
<connection>
<GID>1529</GID>
<name>IN_0</name></connection>
<intersection>718.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>1709</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>717.5,1429.5,719,1429.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_1</name></connection>
<intersection>717.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>717.5,1423,717.5,1429.5</points>
<intersection>1423 21</intersection>
<intersection>1429.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712.5,1423,717.5,1423</points>
<connection>
<GID>1530</GID>
<name>IN_0</name></connection>
<intersection>717.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>1710</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>712.5,1425.5,716.5,1425.5</points>
<connection>
<GID>1531</GID>
<name>IN_0</name></connection>
<intersection>716.5 23</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>716.5,1425.5,716.5,1430.5</points>
<intersection>1425.5 15</intersection>
<intersection>1430.5 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>716.5,1430.5,719,1430.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_2</name></connection>
<intersection>716.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>1711</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>715.5,1431.5,719,1431.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_3</name></connection>
<intersection>715.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>715.5,1428,715.5,1431.5</points>
<intersection>1428 21</intersection>
<intersection>1431.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712.5,1428,715.5,1428</points>
<connection>
<GID>1532</GID>
<name>IN_0</name></connection>
<intersection>715.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>1712</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>714.5,1432.5,719,1432.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_4</name></connection>
<intersection>714.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>714.5,1430.5,714.5,1432.5</points>
<intersection>1430.5 21</intersection>
<intersection>1432.5 15</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712.5,1430.5,714.5,1430.5</points>
<connection>
<GID>1533</GID>
<name>IN_0</name></connection>
<intersection>714.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>1713</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>714,1433.5,719,1433.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_5</name></connection>
<intersection>714 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>714,1432.5,714,1433.5</points>
<intersection>1432.5 21</intersection>
<intersection>1433.5 1</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712.5,1432.5,714,1432.5</points>
<connection>
<GID>1535</GID>
<name>IN_0</name></connection>
<intersection>714 20</intersection></hsegment></shape></wire>
<wire>
<ID>1714</ID>
<shape>
<hsegment>
<ID>15</ID>
<points>714,1434.5,719,1434.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_6</name></connection>
<intersection>714 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>714,1434.5,714,1435</points>
<intersection>1434.5 15</intersection>
<intersection>1435 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>712,1435,714,1435</points>
<connection>
<GID>1534</GID>
<name>IN_0</name></connection>
<intersection>714 20</intersection></hsegment></shape></wire>
<wire>
<ID>1715</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>712,1437.5,715,1437.5</points>
<connection>
<GID>1536</GID>
<name>IN_0</name></connection>
<intersection>715 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>715,1435.5,715,1437.5</points>
<intersection>1435.5 25</intersection>
<intersection>1437.5 1</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>715,1435.5,719,1435.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_7</name></connection>
<intersection>715 24</intersection></hsegment></shape></wire>
<wire>
<ID>1716</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>755.5,1438.5,761.5,1438.5</points>
<connection>
<GID>1537</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1541</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1717</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>755.5,1437.5,756.5,1437.5</points>
<connection>
<GID>1537</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1540</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1718</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>755.5,1436.5,761.5,1436.5</points>
<connection>
<GID>1537</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1539</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1719</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>755.5,1435.5,756.5,1435.5</points>
<connection>
<GID>1537</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1538</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>751.5,1441.5,751.5,1444.5</points>
<connection>
<GID>1537</GID>
<name>count_enable</name></connection>
<connection>
<GID>1542</GID>
<name>OUT</name></connection>
<intersection>1442 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>739.5,1442,751.5,1442</points>
<intersection>739.5 5</intersection>
<intersection>751.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>739.5,1432.5,739.5,1442</points>
<intersection>1432.5 6</intersection>
<intersection>1442 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>739.5,1432.5,741,1432.5</points>
<connection>
<GID>1548</GID>
<name>IN_0</name></connection>
<intersection>739.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>1721</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>753.5,1450.5,753.5,1452.5</points>
<connection>
<GID>1542</GID>
<name>IN_0</name></connection>
<connection>
<GID>1543</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>751.5,1450.5,751.5,1452.5</points>
<connection>
<GID>1542</GID>
<name>IN_1</name></connection>
<connection>
<GID>1544</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>749.5,1450.5,749.5,1452.5</points>
<connection>
<GID>1542</GID>
<name>IN_2</name></connection>
<connection>
<GID>1546</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1724</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>750.5,1431.5,750.5,1432.5</points>
<connection>
<GID>1537</GID>
<name>clock</name></connection>
<intersection>1431.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>747,1431.5,750.5,1431.5</points>
<connection>
<GID>1548</GID>
<name>OUT</name></connection>
<intersection>750.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>752.5,1429,752.5,1432.5</points>
<connection>
<GID>1537</GID>
<name>clear</name></connection>
<intersection>1429 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>752.5,1429,758,1429</points>
<connection>
<GID>1556</GID>
<name>OUT</name></connection>
<intersection>752.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1726</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>764,1430,768.5,1430</points>
<connection>
<GID>1556</GID>
<name>IN_1</name></connection>
<intersection>768.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>768.5,1430,768.5,1430.5</points>
<connection>
<GID>1561</GID>
<name>IN_0</name></connection>
<intersection>1430 1</intersection></vsegment></shape></wire>
<wire>
<ID>1727</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>764,1428,765,1428</points>
<connection>
<GID>1556</GID>
<name>IN_0</name></connection>
<intersection>765 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>765,1427.5,765,1428</points>
<connection>
<GID>1563</GID>
<name>IN_0</name></connection>
<intersection>1428 1</intersection></vsegment></shape></wire>
<wire>
<ID>1728</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>556.5,1430,561,1430</points>
<connection>
<GID>1565</GID>
<name>OUT</name></connection>
<connection>
<GID>1567</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>561,1426.5,561,1428</points>
<connection>
<GID>1567</GID>
<name>IN_1</name></connection>
<intersection>1426.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>559,1426.5,561,1426.5</points>
<connection>
<GID>1570</GID>
<name>OUT_0</name></connection>
<intersection>561 0</intersection></hsegment></shape></wire>
<wire>
<ID>1730</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>550.5,1426.5,555,1426.5</points>
<connection>
<GID>1570</GID>
<name>IN_0</name></connection>
<intersection>550.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>550.5,1426.5,550.5,1434.5</points>
<connection>
<GID>1565</GID>
<name>IN_1</name></connection>
<intersection>1426.5 1</intersection>
<intersection>1434.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>530,1434.5,550.5,1434.5</points>
<connection>
<GID>1199</GID>
<name>OUT_0</name></connection>
<intersection>550.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>567.5,1423,567.5,1429</points>
<connection>
<GID>1607</GID>
<name>IN_0</name></connection>
<intersection>1429 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>567,1429,567.5,1429</points>
<connection>
<GID>1567</GID>
<name>OUT</name></connection>
<intersection>567.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1732</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>573.5,1422,575.5,1422</points>
<connection>
<GID>1607</GID>
<name>OUT</name></connection>
<connection>
<GID>1605</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1733</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>565.5,1421,567.5,1421</points>
<connection>
<GID>1609</GID>
<name>OUT</name></connection>
<connection>
<GID>1607</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1734</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>556.5,1422,559.5,1422</points>
<connection>
<GID>1610</GID>
<name>OUT</name></connection>
<connection>
<GID>1609</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1735</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>547,1421,550.5,1421</points>
<connection>
<GID>1613</GID>
<name>IN_0</name></connection>
<connection>
<GID>1610</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1736</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>544.5,1431,550.5,1431</points>
<connection>
<GID>1615</GID>
<name>IN_0</name></connection>
<connection>
<GID>1565</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>558.5,1411.5,558.5,1420</points>
<intersection>1411.5 2</intersection>
<intersection>1420 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>558.5,1420,559.5,1420</points>
<connection>
<GID>1609</GID>
<name>IN_1</name></connection>
<intersection>558.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>553.5,1411.5,558.5,1411.5</points>
<connection>
<GID>1547</GID>
<name>OUT</name></connection>
<intersection>558.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1738</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>545.5,1412.5,547.5,1412.5</points>
<connection>
<GID>1549</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1547</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1739</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>540,1410.5,547.5,1410.5</points>
<connection>
<GID>1552</GID>
<name>IN_0</name></connection>
<connection>
<GID>1547</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>717.5,1436.5,717.5,1444.5</points>
<connection>
<GID>1612</GID>
<name>OUT_0</name></connection>
<intersection>1436.5 111</intersection>
<intersection>1437.5 112</intersection>
<intersection>1438.5 105</intersection>
<intersection>1439.5 106</intersection>
<intersection>1440.5 107</intersection>
<intersection>1441.5 108</intersection>
<intersection>1442.5 109</intersection>
<intersection>1443.5 110</intersection></vsegment>
<hsegment>
<ID>105</ID>
<points>717.5,1438.5,719,1438.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_10</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>106</ID>
<points>717.5,1439.5,719,1439.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_11</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>107</ID>
<points>717.5,1440.5,719,1440.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_12</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>108</ID>
<points>717.5,1441.5,719,1441.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_13</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>109</ID>
<points>717.5,1442.5,719,1442.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_14</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>110</ID>
<points>717.5,1443.5,719,1443.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_15</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>111</ID>
<points>717.5,1436.5,719,1436.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_8</name></connection>
<intersection>717.5 0</intersection></hsegment>
<hsegment>
<ID>112</ID>
<points>717.5,1437.5,719,1437.5</points>
<connection>
<GID>1524</GID>
<name>ADDRESS_9</name></connection>
<intersection>717.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1741</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>738,1435.5,738,1438</points>
<connection>
<GID>1614</GID>
<name>OUT_0</name></connection>
<intersection>1435.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>737,1435.5,738,1435.5</points>
<connection>
<GID>1524</GID>
<name>ENABLE_0</name></connection>
<intersection>738 0</intersection></hsegment></shape></wire>
<wire>
<ID>1742</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557.5,1506,559,1506</points>
<connection>
<GID>1484</GID>
<name>OUT_0</name></connection>
<intersection>559 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>559,1497,559,1506</points>
<intersection>1497 3</intersection>
<intersection>1506 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>559,1497,577,1497</points>
<connection>
<GID>1490</GID>
<name>IN_0</name></connection>
<intersection>559 2</intersection></hsegment></shape></wire>
<wire>
<ID>1743</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>740.5,1423,740.5,1430.5</points>
<intersection>1423 2</intersection>
<intersection>1430.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>740.5,1430.5,741,1430.5</points>
<connection>
<GID>1548</GID>
<name>IN_1</name></connection>
<intersection>740.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>740.5,1423,742.5,1423</points>
<connection>
<GID>1611</GID>
<name>OUT</name></connection>
<intersection>740.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1744</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>748.5,1424,750.5,1424</points>
<connection>
<GID>1611</GID>
<name>IN_1</name></connection>
<connection>
<GID>1553</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1745</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>748.5,1422,753,1422</points>
<connection>
<GID>1611</GID>
<name>IN_0</name></connection>
<connection>
<GID>1551</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1746</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1457,562.5,1457</points>
<connection>
<GID>1275</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1747</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1455,562.5,1455</points>
<connection>
<GID>1276</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1748</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1453,562.5,1453</points>
<connection>
<GID>1277</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1749</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1451,562.5,1451</points>
<connection>
<GID>1278</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1750</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1449,562.5,1449</points>
<connection>
<GID>1279</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1751</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>562,1447,562.5,1447</points>
<connection>
<GID>1280</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1752</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>561.5,1445,562.5,1445</points>
<connection>
<GID>1283</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1753</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>561,1443,562.5,1443</points>
<connection>
<GID>1284</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1754</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1448,562.5,1448</points>
<connection>
<GID>1309</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1755</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1446,562.5,1446</points>
<connection>
<GID>1310</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1756</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1444,562.5,1444</points>
<connection>
<GID>1285</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1757</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1442,562.5,1442</points>
<connection>
<GID>1286</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1758</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1456,562.5,1456</points>
<connection>
<GID>1287</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1759</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1454,562.5,1454</points>
<connection>
<GID>1289</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1760</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1452,562.5,1452</points>
<connection>
<GID>1290</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1761</ID>
<shape>
<hsegment>
<ID>8</ID>
<points>553.5,1450,562.5,1450</points>
<connection>
<GID>1307</GID>
<name>IN_0</name></connection>
<connection>
<GID>1621</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1762</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1442,590.5,1442</points>
<connection>
<GID>1621</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1261</GID>
<name>IN_0</name></connection>
<intersection>578 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>578,1442,578,1463</points>
<intersection>1442 1</intersection>
<intersection>1463 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1463,578,1463</points>
<connection>
<GID>1620</GID>
<name>OUT_0</name></connection>
<intersection>578 7</intersection></hsegment></shape></wire>
<wire>
<ID>1763</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1443,590.5,1443</points>
<connection>
<GID>1621</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1261</GID>
<name>IN_1</name></connection>
<intersection>578.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>578.5,1443,578.5,1464</points>
<intersection>1443 1</intersection>
<intersection>1464 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1464,578.5,1464</points>
<connection>
<GID>1620</GID>
<name>OUT_1</name></connection>
<intersection>578.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1764</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1444,590.5,1444</points>
<connection>
<GID>1621</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1261</GID>
<name>IN_2</name></connection>
<intersection>579 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>579,1444,579,1465</points>
<intersection>1444 1</intersection>
<intersection>1465 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1465,579,1465</points>
<connection>
<GID>1620</GID>
<name>OUT_2</name></connection>
<intersection>579 7</intersection></hsegment></shape></wire>
<wire>
<ID>1765</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1445,590.5,1445</points>
<connection>
<GID>1621</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1261</GID>
<name>IN_3</name></connection>
<intersection>579.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>579.5,1445,579.5,1466</points>
<intersection>1445 1</intersection>
<intersection>1466 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1466,579.5,1466</points>
<connection>
<GID>1620</GID>
<name>OUT_3</name></connection>
<intersection>579.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1766</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1446,590.5,1446</points>
<connection>
<GID>1621</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1261</GID>
<name>IN_4</name></connection>
<intersection>580 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>580,1446,580,1467</points>
<intersection>1446 1</intersection>
<intersection>1467 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1467,580,1467</points>
<connection>
<GID>1620</GID>
<name>OUT_4</name></connection>
<intersection>580 7</intersection></hsegment></shape></wire>
<wire>
<ID>1767</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1447,590.5,1447</points>
<connection>
<GID>1621</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1261</GID>
<name>IN_5</name></connection>
<intersection>580.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>580.5,1447,580.5,1468</points>
<intersection>1447 1</intersection>
<intersection>1468 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>577.5,1468,580.5,1468</points>
<connection>
<GID>1620</GID>
<name>OUT_5</name></connection>
<intersection>580.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1768</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1448,590.5,1448</points>
<connection>
<GID>1621</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1261</GID>
<name>IN_6</name></connection>
<intersection>581 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>581,1448,581,1469</points>
<intersection>1448 1</intersection>
<intersection>1469 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1469,581,1469</points>
<connection>
<GID>1620</GID>
<name>OUT_6</name></connection>
<intersection>581 7</intersection></hsegment></shape></wire>
<wire>
<ID>1769</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1449,590.5,1449</points>
<connection>
<GID>1621</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1261</GID>
<name>IN_7</name></connection>
<intersection>581.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>581.5,1449,581.5,1470</points>
<intersection>1449 1</intersection>
<intersection>1470 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1470,581.5,1470</points>
<connection>
<GID>1620</GID>
<name>OUT_7</name></connection>
<intersection>581.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1770</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1450,590.5,1450</points>
<connection>
<GID>1621</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1261</GID>
<name>IN_8</name></connection>
<intersection>582 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>582,1450,582,1471</points>
<intersection>1450 1</intersection>
<intersection>1471 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1471,582,1471</points>
<connection>
<GID>1620</GID>
<name>OUT_8</name></connection>
<intersection>582 7</intersection></hsegment></shape></wire>
<wire>
<ID>1771</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1451,590.5,1451</points>
<connection>
<GID>1621</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1261</GID>
<name>IN_9</name></connection>
<intersection>582.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>582.5,1451,582.5,1472</points>
<intersection>1451 1</intersection>
<intersection>1472 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1472,582.5,1472</points>
<connection>
<GID>1620</GID>
<name>OUT_9</name></connection>
<intersection>582.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1772</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1452,590.5,1452</points>
<connection>
<GID>1621</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1261</GID>
<name>IN_10</name></connection>
<intersection>583 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>583,1452,583,1473</points>
<intersection>1452 1</intersection>
<intersection>1473 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1473,583,1473</points>
<connection>
<GID>1620</GID>
<name>OUT_10</name></connection>
<intersection>583 7</intersection></hsegment></shape></wire>
<wire>
<ID>1773</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1453,590.5,1453</points>
<connection>
<GID>1621</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1261</GID>
<name>IN_11</name></connection>
<intersection>583.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>583.5,1453,583.5,1474</points>
<intersection>1453 1</intersection>
<intersection>1474 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1474,583.5,1474</points>
<connection>
<GID>1620</GID>
<name>OUT_11</name></connection>
<intersection>583.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1774</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1454,590.5,1454</points>
<connection>
<GID>1621</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1261</GID>
<name>IN_12</name></connection>
<intersection>584 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>584,1454,584,1475</points>
<intersection>1454 1</intersection>
<intersection>1475 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1475,584,1475</points>
<connection>
<GID>1620</GID>
<name>OUT_12</name></connection>
<intersection>584 7</intersection></hsegment></shape></wire>
<wire>
<ID>1775</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1455,590.5,1455</points>
<connection>
<GID>1621</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1261</GID>
<name>IN_13</name></connection>
<intersection>584.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>584.5,1455,584.5,1476</points>
<intersection>1455 1</intersection>
<intersection>1476 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1476,584.5,1476</points>
<connection>
<GID>1620</GID>
<name>OUT_13</name></connection>
<intersection>584.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1776</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1456,590.5,1456</points>
<connection>
<GID>1621</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1261</GID>
<name>IN_14</name></connection>
<intersection>585 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>585,1456,585,1477</points>
<intersection>1456 1</intersection>
<intersection>1477 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1477,585,1477</points>
<connection>
<GID>1620</GID>
<name>OUT_14</name></connection>
<intersection>585 7</intersection></hsegment></shape></wire>
<wire>
<ID>1777</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>566.5,1457,590.5,1457</points>
<connection>
<GID>1621</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1261</GID>
<name>IN_15</name></connection>
<intersection>585.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>585.5,1457,585.5,1478</points>
<intersection>1457 1</intersection>
<intersection>1478 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>577.5,1478,585.5,1478</points>
<connection>
<GID>1620</GID>
<name>OUT_15</name></connection>
<intersection>585.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>1778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,1458.5,564.5,1460.5</points>
<connection>
<GID>1621</GID>
<name>ENABLE_0</name></connection>
<intersection>1460.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>561,1460.5,564.5,1460.5</points>
<connection>
<GID>1622</GID>
<name>OUT_0</name></connection>
<intersection>564.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1321</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1483,632,1483</points>
<connection>
<GID>1195</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1312</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1322</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1481,632,1481</points>
<connection>
<GID>1195</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1313</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1479,632,1479</points>
<connection>
<GID>1195</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1314</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1324</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1477,632,1477</points>
<connection>
<GID>1195</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1315</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1325</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1475,632,1475</points>
<connection>
<GID>1195</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1316</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1326</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1473,632,1473</points>
<connection>
<GID>1195</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1317</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1327</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1471,632,1471</points>
<connection>
<GID>1195</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1318</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1469,632,1469</points>
<connection>
<GID>1195</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1319</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1329</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1482,625,1482</points>
<connection>
<GID>1195</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1320</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1480,625,1480</points>
<connection>
<GID>1195</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1321</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1331</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1478,625,1478</points>
<connection>
<GID>1195</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1322</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1332</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1476,625,1476</points>
<connection>
<GID>1195</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1323</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1333</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1474,625,1474</points>
<connection>
<GID>1195</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1324</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1334</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1472,625,1472</points>
<connection>
<GID>1195</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1325</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1335</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1470,625,1470</points>
<connection>
<GID>1195</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1326</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1336</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1468,625,1468</points>
<connection>
<GID>1195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1327</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534.5,1474,534.5,1490.5</points>
<intersection>1474 2</intersection>
<intersection>1490.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>534.5,1490.5,536,1490.5</points>
<connection>
<GID>1196</GID>
<name>N_in0</name></connection>
<intersection>534.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525,1474,534.5,1474</points>
<connection>
<GID>1197</GID>
<name>OUT_8</name></connection>
<intersection>534.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1338</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>538,1490.5,539,1490.5</points>
<connection>
<GID>1196</GID>
<name>N_in1</name></connection>
<connection>
<GID>1243</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>532.5,1462.5,532.5,1466</points>
<intersection>1462.5 2</intersection>
<intersection>1466 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1466,532.5,1466</points>
<connection>
<GID>1197</GID>
<name>OUT_0</name></connection>
<intersection>532.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>532.5,1462.5,540,1462.5</points>
<connection>
<GID>1271</GID>
<name>IN_0</name></connection>
<intersection>532.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,1466,539,1467</points>
<intersection>1466 2</intersection>
<intersection>1467 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1467,539,1467</points>
<connection>
<GID>1197</GID>
<name>OUT_1</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,1466,540,1466</points>
<connection>
<GID>1200</GID>
<name>IN_0</name></connection>
<intersection>539 0</intersection></hsegment></shape></wire>
<wire>
<ID>1341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>575.5,1479.5,575.5,1484</points>
<connection>
<GID>1620</GID>
<name>ENABLE_0</name></connection>
<intersection>1484 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>574,1484,575.5,1484</points>
<connection>
<GID>1288</GID>
<name>IN_0</name></connection>
<intersection>575.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1342</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1496,699.5,1496</points>
<connection>
<GID>1281</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1343</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1494,699.5,1494</points>
<connection>
<GID>1281</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1213</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1492,699.5,1492</points>
<connection>
<GID>1281</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1215</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1490,699.5,1490</points>
<connection>
<GID>1281</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1217</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1488,699.5,1488</points>
<connection>
<GID>1281</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1244</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>539,1468,539,1469</points>
<intersection>1468 1</intersection>
<intersection>1469 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1468,539,1468</points>
<connection>
<GID>1197</GID>
<name>OUT_2</name></connection>
<intersection>539 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>539,1469,540,1469</points>
<connection>
<GID>1201</GID>
<name>IN_0</name></connection>
<intersection>539 0</intersection></hsegment></shape></wire>
<wire>
<ID>1348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1486,699.5,1486</points>
<connection>
<GID>1281</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1245</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>538,1469,538,1472</points>
<intersection>1469 1</intersection>
<intersection>1472 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1469,538,1469</points>
<connection>
<GID>1197</GID>
<name>OUT_3</name></connection>
<intersection>538 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>538,1472,540,1472</points>
<connection>
<GID>1218</GID>
<name>IN_0</name></connection>
<intersection>538 0</intersection></hsegment></shape></wire>
<wire>
<ID>1350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1484,699.5,1484</points>
<connection>
<GID>1281</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1246</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1351</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535.5,1471,535.5,1481</points>
<intersection>1471 2</intersection>
<intersection>1481 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535.5,1481,540,1481</points>
<connection>
<GID>1241</GID>
<name>IN_0</name></connection>
<intersection>535.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525,1471,535.5,1471</points>
<connection>
<GID>1197</GID>
<name>OUT_5</name></connection>
<intersection>535.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>535,1472,535,1484</points>
<intersection>1472 2</intersection>
<intersection>1484 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>535,1484,540,1484</points>
<connection>
<GID>1242</GID>
<name>IN_0</name></connection>
<intersection>535 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525,1472,535,1472</points>
<connection>
<GID>1197</GID>
<name>OUT_6</name></connection>
<intersection>535 0</intersection></hsegment></shape></wire>
<wire>
<ID>1353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>515.5,1481,519,1481</points>
<connection>
<GID>1250</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1197</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>1354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,1469,517,1472</points>
<intersection>1469 1</intersection>
<intersection>1472 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,1469,519,1469</points>
<connection>
<GID>1197</GID>
<name>IN_3</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,1472,517,1472</points>
<connection>
<GID>1251</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment></shape></wire>
<wire>
<ID>1355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,1468,516.5,1469</points>
<intersection>1468 1</intersection>
<intersection>1469 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516.5,1468,519,1468</points>
<connection>
<GID>1197</GID>
<name>IN_2</name></connection>
<intersection>516.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,1469,516.5,1469</points>
<connection>
<GID>1253</GID>
<name>IN_0</name></connection>
<intersection>516.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>516.5,1466,516.5,1467</points>
<intersection>1466 2</intersection>
<intersection>1467 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>516.5,1467,519,1467</points>
<connection>
<GID>1197</GID>
<name>IN_1</name></connection>
<intersection>516.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,1466,516.5,1466</points>
<connection>
<GID>1254</GID>
<name>IN_0</name></connection>
<intersection>516.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>517,1463,517,1466</points>
<intersection>1463 2</intersection>
<intersection>1466 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>517,1466,519,1466</points>
<connection>
<GID>1197</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>514,1463,517,1463</points>
<connection>
<GID>1255</GID>
<name>IN_0</name></connection>
<intersection>517 0</intersection></hsegment></shape></wire>
<wire>
<ID>1358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>534,1475,534,1493</points>
<intersection>1475 1</intersection>
<intersection>1493 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1475,534,1475</points>
<connection>
<GID>1197</GID>
<name>OUT_9</name></connection>
<intersection>534 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>534,1493,539,1493</points>
<connection>
<GID>1249</GID>
<name>IN_0</name></connection>
<intersection>534 0</intersection></hsegment></shape></wire>
<wire>
<ID>1359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>680,1406.5,680,1434</points>
<intersection>1406.5 1</intersection>
<intersection>1428 3</intersection>
<intersection>1434 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>677.5,1406.5,680,1406.5</points>
<connection>
<GID>1571</GID>
<name>ENABLE_0</name></connection>
<intersection>680 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>680,1434,686,1434</points>
<connection>
<GID>1252</GID>
<name>IN_0</name></connection>
<intersection>680 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>678,1428,680,1428</points>
<connection>
<GID>1562</GID>
<name>ENABLE_0</name></connection>
<intersection>680 0</intersection></hsegment></shape></wire>
<wire>
<ID>1360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>685,1404,685,1429</points>
<connection>
<GID>1608</GID>
<name>IN_0</name></connection>
<intersection>1406 2</intersection>
<intersection>1429 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>678,1429,685,1429</points>
<connection>
<GID>1562</GID>
<name>write_enable</name></connection>
<intersection>685 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>685,1406,686.5,1406</points>
<connection>
<GID>1572</GID>
<name>ENABLE_0</name></connection>
<intersection>685 0</intersection></hsegment></shape></wire>
<wire>
<ID>1361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>543,1423,543,1425</points>
<intersection>1423 1</intersection>
<intersection>1425 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>543,1423,550.5,1423</points>
<connection>
<GID>1610</GID>
<name>IN_0</name></connection>
<intersection>543 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>535,1425,543,1425</points>
<connection>
<GID>1204</GID>
<name>OUT_0</name></connection>
<intersection>543 0</intersection></hsegment></shape></wire>
<wire>
<ID>1362</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1482,699.5,1482</points>
<connection>
<GID>1281</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1247</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>537,1470,537,1475</points>
<intersection>1470 2</intersection>
<intersection>1475 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>537,1475,540,1475</points>
<connection>
<GID>1239</GID>
<name>IN_0</name></connection>
<intersection>537 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>525,1470,537,1470</points>
<connection>
<GID>1197</GID>
<name>OUT_4</name></connection>
<intersection>537 0</intersection></hsegment></shape></wire>
<wire>
<ID>1364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1497,691,1497</points>
<connection>
<GID>1281</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1248</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1495,691,1495</points>
<connection>
<GID>1281</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1256</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1493,691,1493</points>
<connection>
<GID>1281</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1257</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1491,691,1491</points>
<connection>
<GID>1281</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1258</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1489,691,1489</points>
<connection>
<GID>1281</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1259</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1487,691,1487</points>
<connection>
<GID>1281</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1262</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1485,691,1485</points>
<connection>
<GID>1281</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1264</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>688,1483,691,1483</points>
<connection>
<GID>1281</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1265</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>533,1477,533,1495.5</points>
<intersection>1477 1</intersection>
<intersection>1495.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1477,533,1477</points>
<connection>
<GID>1197</GID>
<name>OUT_11</name></connection>
<intersection>533 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>533,1495.5,541,1495.5</points>
<connection>
<GID>1240</GID>
<name>IN_0</name></connection>
<intersection>533 0</intersection></hsegment></shape></wire>
<wire>
<ID>1373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621,1484.5,621,1488</points>
<connection>
<GID>1195</GID>
<name>ENABLE_0</name></connection>
<intersection>1488 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>621,1488,639,1488</points>
<connection>
<GID>1202</GID>
<name>OUT</name></connection>
<intersection>621 0</intersection></hsegment></shape></wire>
<wire>
<ID>1374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557.5,1514.5,563,1514.5</points>
<connection>
<GID>1269</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1266</GID>
<name>IN_0</name></connection>
<intersection>561 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>561,1508,561,1514.5</points>
<connection>
<GID>1268</GID>
<name>IN_0</name></connection>
<intersection>1514.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>647.5,1489,647.5,1489.5</points>
<intersection>1489 1</intersection>
<intersection>1489.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,1489,647.5,1489</points>
<connection>
<GID>1202</GID>
<name>IN_2</name></connection>
<intersection>647.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>647.5,1489.5,649,1489.5</points>
<connection>
<GID>1308</GID>
<name>IN_0</name></connection>
<intersection>647.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1376</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>646,1487,649.5,1487</points>
<connection>
<GID>1202</GID>
<name>IN_1</name></connection>
<connection>
<GID>1198</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>647.5,1484.5,647.5,1485</points>
<intersection>1484.5 2</intersection>
<intersection>1485 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,1485,647.5,1485</points>
<connection>
<GID>1202</GID>
<name>IN_0</name></connection>
<intersection>647.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>647.5,1484.5,649.5,1484.5</points>
<connection>
<GID>1205</GID>
<name>IN_0</name></connection>
<intersection>647.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>686,1498.5,686,1501</points>
<connection>
<GID>1281</GID>
<name>ENABLE_0</name></connection>
<intersection>1501 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>686,1501,694,1501</points>
<connection>
<GID>1282</GID>
<name>IN_0</name></connection>
<intersection>686 0</intersection></hsegment></shape></wire>
<wire>
<ID>1379</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1467,573.5,1467</points>
<connection>
<GID>1293</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1380</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1463,573.5,1463</points>
<connection>
<GID>1291</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1465,573.5,1465</points>
<connection>
<GID>1292</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1382</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1469,573.5,1469</points>
<connection>
<GID>1294</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1383</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1471,573.5,1471</points>
<connection>
<GID>1295</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1384</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1473,573.5,1473</points>
<connection>
<GID>1296</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1385</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1475,573.5,1475</points>
<connection>
<GID>1297</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1386</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>567.5,1477,573.5,1477</points>
<connection>
<GID>1298</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1387</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,1464,573.5,1464</points>
<connection>
<GID>1299</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1388</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,1478,573.5,1478</points>
<connection>
<GID>1306</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1620</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1389</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>532,1516.5,577,1516.5</points>
<intersection>532 5</intersection>
<intersection>562.5 6</intersection>
<intersection>577 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>577,1507.5,577,1516.5</points>
<intersection>1507.5 4</intersection>
<intersection>1516.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>577,1507.5,578.5,1507.5</points>
<connection>
<GID>1208</GID>
<name>IN_0</name></connection>
<intersection>577 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>532,1506.5,532,1516.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>1516.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>562.5,1516.5,562.5,1518.5</points>
<intersection>1516.5 1</intersection>
<intersection>1518.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>557.5,1518.5,562.5,1518.5</points>
<connection>
<GID>1209</GID>
<name>OUT_0</name></connection>
<intersection>562.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>1390</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>559,1510.5,559,1512.5</points>
<intersection>1510.5 4</intersection>
<intersection>1512.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>559,1512.5,563,1512.5</points>
<connection>
<GID>1266</GID>
<name>IN_1</name></connection>
<intersection>559 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>558.5,1510.5,559,1510.5</points>
<connection>
<GID>1219</GID>
<name>OUT_0</name></connection>
<intersection>559 0</intersection></hsegment></shape></wire>
<wire>
<ID>1391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531,1479,531,1499</points>
<intersection>1479 1</intersection>
<intersection>1499 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>525,1479,531,1479</points>
<connection>
<GID>1197</GID>
<name>OUT_13</name></connection>
<intersection>531 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>531,1499,541,1499</points>
<connection>
<GID>1222</GID>
<name>IN_0</name></connection>
<intersection>531 0</intersection></hsegment></shape></wire>
<wire>
<ID>1392</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>532,1498,578.5,1498</points>
<intersection>532 2</intersection>
<intersection>577 3</intersection>
<intersection>578.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>532,1498,532,1504.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>1498 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>577,1498,577,1505.5</points>
<connection>
<GID>1270</GID>
<name>OUT</name></connection>
<intersection>1498 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>578.5,1498,578.5,1505.5</points>
<connection>
<GID>1208</GID>
<name>IN_1</name></connection>
<intersection>1498 1</intersection></vsegment></shape></wire>
<wire>
<ID>1393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>570,1506.5,570,1513.5</points>
<intersection>1506.5 1</intersection>
<intersection>1513.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>570,1506.5,571,1506.5</points>
<connection>
<GID>1270</GID>
<name>IN_0</name></connection>
<intersection>570 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>569,1513.5,570,1513.5</points>
<connection>
<GID>1266</GID>
<name>OUT</name></connection>
<intersection>570 0</intersection></hsegment></shape></wire>
<wire>
<ID>1394</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>653,1497,656,1497</points>
<connection>
<GID>1220</GID>
<name>IN_1</name></connection>
<intersection>656 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>656,1496.5,656,1497</points>
<intersection>1496.5 5</intersection>
<intersection>1497 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>656,1496.5,657.5,1496.5</points>
<connection>
<GID>1203</GID>
<name>IN_0</name></connection>
<intersection>656 4</intersection></hsegment></shape></wire>
<wire>
<ID>1395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>654.5,1493,654.5,1495</points>
<intersection>1493 3</intersection>
<intersection>1495 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653,1495,654.5,1495</points>
<connection>
<GID>1220</GID>
<name>IN_0</name></connection>
<intersection>654.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>654.5,1493,655,1493</points>
<connection>
<GID>1221</GID>
<name>IN_0</name></connection>
<intersection>654.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>646.5,1491,646.5,1496</points>
<intersection>1491 1</intersection>
<intersection>1496 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>646,1491,646.5,1491</points>
<connection>
<GID>1202</GID>
<name>IN_3</name></connection>
<intersection>646.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>646.5,1496,647,1496</points>
<connection>
<GID>1220</GID>
<name>OUT</name></connection>
<intersection>646.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1397</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557,1500.5,562.5,1500.5</points>
<connection>
<GID>1206</GID>
<name>CLK</name></connection>
<connection>
<GID>1267</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>561,1502.5,561,1504</points>
<connection>
<GID>1268</GID>
<name>OUT_0</name></connection>
<intersection>1502.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>561,1502.5,562.5,1502.5</points>
<connection>
<GID>1267</GID>
<name>IN_0</name></connection>
<intersection>561 0</intersection></hsegment></shape></wire>
<wire>
<ID>1399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>569.5,1501.5,569.5,1504.5</points>
<intersection>1501.5 2</intersection>
<intersection>1504.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>569.5,1504.5,571,1504.5</points>
<connection>
<GID>1270</GID>
<name>IN_1</name></connection>
<intersection>569.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>568.5,1501.5,569.5,1501.5</points>
<connection>
<GID>1267</GID>
<name>OUT</name></connection>
<intersection>569.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1400</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1422,645.5,1422</points>
<connection>
<GID>1328</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1401</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1424,645.5,1424</points>
<connection>
<GID>1311</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1402</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1436,645.5,1436</points>
<connection>
<GID>1357</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1403</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1434,645.5,1434</points>
<connection>
<GID>1359</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1404</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1432,645.5,1432</points>
<connection>
<GID>1361</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1405</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1430,645.5,1430</points>
<connection>
<GID>1363</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1406</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1428,645.5,1428</points>
<connection>
<GID>1364</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1407</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>644.5,1426,645.5,1426</points>
<connection>
<GID>1365</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1408</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1423,645.5,1423</points>
<connection>
<GID>1329</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1409</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1421,645.5,1421</points>
<connection>
<GID>1330</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1410</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1435,645.5,1435</points>
<connection>
<GID>1331</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1411</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1433,645.5,1433</points>
<connection>
<GID>1332</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1412</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1431,645.5,1431</points>
<connection>
<GID>1334</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1413</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1429,645.5,1429</points>
<connection>
<GID>1352</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1427,645.5,1427</points>
<connection>
<GID>1353</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>638,1425,645.5,1425</points>
<connection>
<GID>1355</GID>
<name>IN_0</name></connection>
<connection>
<GID>1564</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1416</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1404,594,1404</points>
<connection>
<GID>1384</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1451,619,1451</points>
<connection>
<GID>1261</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1333</GID>
<name>IN_9</name></connection>
<intersection>607 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>607,1451,607,1500</points>
<intersection>1451 1</intersection>
<intersection>1477 13</intersection>
<intersection>1500 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>607,1477,619,1477</points>
<connection>
<GID>1195</GID>
<name>IN_9</name></connection>
<intersection>607 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>607,1500,633,1500</points>
<connection>
<GID>1226</GID>
<name>IN_0</name></connection>
<intersection>607 12</intersection></hsegment></shape></wire>
<wire>
<ID>1418</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1457,619,1457</points>
<connection>
<GID>1261</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1333</GID>
<name>IN_15</name></connection>
<intersection>601 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>601,1457,601,1506</points>
<intersection>1457 1</intersection>
<intersection>1483 13</intersection>
<intersection>1506 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>601,1483,619,1483</points>
<connection>
<GID>1195</GID>
<name>IN_15</name></connection>
<intersection>601 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>601,1506,633,1506</points>
<connection>
<GID>1223</GID>
<name>IN_0</name></connection>
<intersection>601 12</intersection></hsegment></shape></wire>
<wire>
<ID>1419</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1455,619,1455</points>
<connection>
<GID>1261</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1333</GID>
<name>IN_13</name></connection>
<intersection>603 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>603,1455,603,1504</points>
<intersection>1455 1</intersection>
<intersection>1481 13</intersection>
<intersection>1504 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>603,1481,619,1481</points>
<connection>
<GID>1195</GID>
<name>IN_13</name></connection>
<intersection>603 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>603,1504,633,1504</points>
<connection>
<GID>1224</GID>
<name>IN_0</name></connection>
<intersection>603 12</intersection></hsegment></shape></wire>
<wire>
<ID>1420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1453,619,1453</points>
<connection>
<GID>1261</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1333</GID>
<name>IN_11</name></connection>
<intersection>605 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>605,1453,605,1502</points>
<intersection>1453 1</intersection>
<intersection>1479 13</intersection>
<intersection>1502 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>605,1479,619,1479</points>
<connection>
<GID>1195</GID>
<name>IN_11</name></connection>
<intersection>605 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>605,1502,633,1502</points>
<connection>
<GID>1225</GID>
<name>IN_0</name></connection>
<intersection>605 12</intersection></hsegment></shape></wire>
<wire>
<ID>1421</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1449,619,1449</points>
<connection>
<GID>1261</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1333</GID>
<name>IN_7</name></connection>
<intersection>609 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>609,1449,609,1498</points>
<intersection>1449 1</intersection>
<intersection>1475 13</intersection>
<intersection>1498 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>609,1475,619,1475</points>
<connection>
<GID>1195</GID>
<name>IN_7</name></connection>
<intersection>609 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>609,1498,633,1498</points>
<connection>
<GID>1227</GID>
<name>IN_0</name></connection>
<intersection>609 12</intersection></hsegment></shape></wire>
<wire>
<ID>1422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1447,619,1447</points>
<connection>
<GID>1261</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1333</GID>
<name>IN_5</name></connection>
<intersection>611 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>611,1447,611,1496</points>
<intersection>1447 1</intersection>
<intersection>1473 13</intersection>
<intersection>1496 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>611,1473,619,1473</points>
<connection>
<GID>1195</GID>
<name>IN_5</name></connection>
<intersection>611 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>611,1496,633,1496</points>
<connection>
<GID>1228</GID>
<name>IN_0</name></connection>
<intersection>611 12</intersection></hsegment></shape></wire>
<wire>
<ID>1423</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1445,619,1445</points>
<connection>
<GID>1261</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1333</GID>
<name>IN_3</name></connection>
<intersection>613 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>613,1445,613,1494</points>
<intersection>1445 1</intersection>
<intersection>1471 13</intersection>
<intersection>1494 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>613,1471,619,1471</points>
<connection>
<GID>1195</GID>
<name>IN_3</name></connection>
<intersection>613 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>613,1494,633,1494</points>
<connection>
<GID>1229</GID>
<name>IN_0</name></connection>
<intersection>613 12</intersection></hsegment></shape></wire>
<wire>
<ID>1424</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,1443,619,1443</points>
<connection>
<GID>1261</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1333</GID>
<name>IN_1</name></connection>
<intersection>615 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>615,1443,615,1492</points>
<intersection>1443 1</intersection>
<intersection>1469 13</intersection>
<intersection>1492 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>615,1469,619,1469</points>
<connection>
<GID>1195</GID>
<name>IN_1</name></connection>
<intersection>615 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>615,1492,633,1492</points>
<connection>
<GID>1230</GID>
<name>IN_0</name></connection>
<intersection>615 12</intersection></hsegment></shape></wire>
<wire>
<ID>1425</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1456,619,1456</points>
<connection>
<GID>1261</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1333</GID>
<name>IN_14</name></connection>
<intersection>602 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>602,1456,602,1505</points>
<intersection>1456 0</intersection>
<intersection>1482 13</intersection>
<intersection>1505 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>602,1482,619,1482</points>
<connection>
<GID>1195</GID>
<name>IN_14</name></connection>
<intersection>602 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>602,1505,626,1505</points>
<connection>
<GID>1231</GID>
<name>IN_0</name></connection>
<intersection>602 12</intersection></hsegment></shape></wire>
<wire>
<ID>1426</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1454,619,1454</points>
<connection>
<GID>1261</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1333</GID>
<name>IN_12</name></connection>
<intersection>604 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>604,1454,604,1503</points>
<intersection>1454 0</intersection>
<intersection>1480 13</intersection>
<intersection>1503 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>604,1480,619,1480</points>
<connection>
<GID>1195</GID>
<name>IN_12</name></connection>
<intersection>604 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>604,1503,626,1503</points>
<connection>
<GID>1232</GID>
<name>IN_0</name></connection>
<intersection>604 12</intersection></hsegment></shape></wire>
<wire>
<ID>1427</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1452,619,1452</points>
<connection>
<GID>1261</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1333</GID>
<name>IN_10</name></connection>
<intersection>606 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>606,1452,606,1501</points>
<intersection>1452 0</intersection>
<intersection>1478 12</intersection>
<intersection>1501 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>606,1478,619,1478</points>
<connection>
<GID>1195</GID>
<name>IN_10</name></connection>
<intersection>606 11</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>606,1501,626,1501</points>
<connection>
<GID>1233</GID>
<name>IN_0</name></connection>
<intersection>606 11</intersection></hsegment></shape></wire>
<wire>
<ID>1428</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1450,619,1450</points>
<connection>
<GID>1261</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1333</GID>
<name>IN_8</name></connection>
<intersection>608 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>608,1450,608,1499</points>
<intersection>1450 0</intersection>
<intersection>1476 12</intersection>
<intersection>1499 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>608,1476,619,1476</points>
<connection>
<GID>1195</GID>
<name>IN_8</name></connection>
<intersection>608 11</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>608,1499,626,1499</points>
<connection>
<GID>1234</GID>
<name>IN_0</name></connection>
<intersection>608 11</intersection></hsegment></shape></wire>
<wire>
<ID>1429</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1448,619,1448</points>
<connection>
<GID>1261</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1333</GID>
<name>IN_6</name></connection>
<intersection>610 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>610,1448,610,1497</points>
<intersection>1448 0</intersection>
<intersection>1474 12</intersection>
<intersection>1497 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>610,1474,619,1474</points>
<connection>
<GID>1195</GID>
<name>IN_6</name></connection>
<intersection>610 11</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>610,1497,626,1497</points>
<connection>
<GID>1235</GID>
<name>IN_0</name></connection>
<intersection>610 11</intersection></hsegment></shape></wire>
<wire>
<ID>1430</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1446,619,1446</points>
<connection>
<GID>1261</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1333</GID>
<name>IN_4</name></connection>
<intersection>612 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>612,1446,612,1495</points>
<intersection>1446 0</intersection>
<intersection>1472 12</intersection>
<intersection>1495 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>612,1472,619,1472</points>
<connection>
<GID>1195</GID>
<name>IN_4</name></connection>
<intersection>612 11</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>612,1495,626,1495</points>
<connection>
<GID>1236</GID>
<name>IN_0</name></connection>
<intersection>612 11</intersection></hsegment></shape></wire>
<wire>
<ID>1431</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1444,619,1444</points>
<connection>
<GID>1261</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1333</GID>
<name>IN_2</name></connection>
<intersection>614 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>614,1444,614,1493</points>
<intersection>1444 0</intersection>
<intersection>1470 13</intersection>
<intersection>1493 19</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>614,1470,619,1470</points>
<connection>
<GID>1195</GID>
<name>IN_2</name></connection>
<intersection>614 12</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>614,1493,626,1493</points>
<connection>
<GID>1237</GID>
<name>IN_0</name></connection>
<intersection>614 12</intersection></hsegment></shape></wire>
<wire>
<ID>1432</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>600.5,1442,619,1442</points>
<connection>
<GID>1261</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1333</GID>
<name>IN_0</name></connection>
<intersection>616 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>616,1442,616,1491</points>
<intersection>1442 0</intersection>
<intersection>1468 12</intersection>
<intersection>1491 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>616,1468,619,1468</points>
<connection>
<GID>1195</GID>
<name>IN_0</name></connection>
<intersection>616 11</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>616,1491,626,1491</points>
<connection>
<GID>1238</GID>
<name>IN_0</name></connection>
<intersection>616 11</intersection></hsegment></shape></wire>
<wire>
<ID>1433</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>621,1458.5,621,1460</points>
<connection>
<GID>1333</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>1335</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1434</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1456,625.5,1456</points>
<connection>
<GID>1333</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1344</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1435</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1454,625.5,1454</points>
<connection>
<GID>1333</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1345</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1436</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1452,625.5,1452</points>
<connection>
<GID>1333</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1346</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1437</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1450,625.5,1450</points>
<connection>
<GID>1333</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1347</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1438</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1448,625.5,1448</points>
<connection>
<GID>1333</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1348</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1439</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1446,625.5,1446</points>
<connection>
<GID>1333</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1349</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1440</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1444,625.5,1444</points>
<connection>
<GID>1333</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1350</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1441</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>623,1442,625.5,1442</points>
<connection>
<GID>1333</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1351</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1442</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1447,632.5,1447</points>
<connection>
<GID>1333</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1341</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1443</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1445,632.5,1445</points>
<connection>
<GID>1333</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1342</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1444</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1443,632.5,1443</points>
<connection>
<GID>1333</GID>
<name>OUT_1</name></connection>
<connection>
<GID>1343</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1445</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1449,632.5,1449</points>
<connection>
<GID>1333</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1340</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1446</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1451,632.5,1451</points>
<connection>
<GID>1333</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1339</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1447</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1453,632.5,1453</points>
<connection>
<GID>1333</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1338</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1448</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1455,632.5,1455</points>
<connection>
<GID>1333</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1337</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1449</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>623,1457,632.5,1457</points>
<connection>
<GID>1333</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1336</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594.5,1437,594.5,1440</points>
<connection>
<GID>1261</GID>
<name>clock</name></connection>
<intersection>1437 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>592.5,1437,594.5,1437</points>
<connection>
<GID>1354</GID>
<name>OUT</name></connection>
<intersection>594.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1451</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>596.5,1437,596.5,1440</points>
<connection>
<GID>1261</GID>
<name>clear</name></connection>
<intersection>1437 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>596.5,1437,602,1437</points>
<connection>
<GID>1356</GID>
<name>OUT</name></connection>
<intersection>596.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>581.5,1438,586.5,1438</points>
<connection>
<GID>1358</GID>
<name>IN_0</name></connection>
<connection>
<GID>1354</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>578,1436,586.5,1436</points>
<connection>
<GID>1360</GID>
<name>IN_0</name></connection>
<connection>
<GID>1354</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1454</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>608,1438,613.5,1438</points>
<connection>
<GID>1356</GID>
<name>IN_1</name></connection>
<connection>
<GID>1362</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1455</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>608,1436,608,1436</points>
<connection>
<GID>1356</GID>
<name>IN_0</name></connection>
<connection>
<GID>1377</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1406,594,1406</points>
<connection>
<GID>1383</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1457</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1408,594,1408</points>
<connection>
<GID>1382</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1410,594,1410</points>
<connection>
<GID>1381</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1459</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1412,594,1412</points>
<connection>
<GID>1380</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1414,594,1414</points>
<connection>
<GID>1379</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1461</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1400,594,1400</points>
<connection>
<GID>1369</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>592.5,1402,594,1402</points>
<connection>
<GID>1368</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1463</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1403,594,1403</points>
<connection>
<GID>1378</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1464</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1405,594,1405</points>
<connection>
<GID>1376</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1465</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1407,594,1407</points>
<connection>
<GID>1375</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1466</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1411,594,1411</points>
<connection>
<GID>1373</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1467</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1413,594,1413</points>
<connection>
<GID>1372</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1468</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1399,594,1399</points>
<connection>
<GID>1371</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1469</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1401,594,1401</points>
<connection>
<GID>1370</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1470</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584,1409,594,1409</points>
<connection>
<GID>1374</GID>
<name>IN_0</name></connection>
<connection>
<GID>1526</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1471</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1411,611.5,1411</points>
<connection>
<GID>1527</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1394</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1472</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1413,611.5,1413</points>
<connection>
<GID>1527</GID>
<name>OUT_14</name></connection>
<connection>
<GID>1393</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1473</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1399,611.5,1399</points>
<connection>
<GID>1527</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1400</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1474</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1401,611.5,1401</points>
<connection>
<GID>1527</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1475</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1403,611.5,1403</points>
<connection>
<GID>1527</GID>
<name>OUT_4</name></connection>
<connection>
<GID>1398</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1476</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1405,611.5,1405</points>
<connection>
<GID>1527</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1397</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1477</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1407,611.5,1407</points>
<connection>
<GID>1527</GID>
<name>OUT_8</name></connection>
<connection>
<GID>1396</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1409,611.5,1409</points>
<connection>
<GID>1527</GID>
<name>OUT_10</name></connection>
<connection>
<GID>1395</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1406,619,1406</points>
<connection>
<GID>1527</GID>
<name>OUT_7</name></connection>
<connection>
<GID>1389</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1480</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1408,619,1408</points>
<connection>
<GID>1527</GID>
<name>OUT_9</name></connection>
<connection>
<GID>1388</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1481</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1410,619,1410</points>
<connection>
<GID>1527</GID>
<name>OUT_11</name></connection>
<connection>
<GID>1387</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1482</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1412,619,1412</points>
<connection>
<GID>1527</GID>
<name>OUT_13</name></connection>
<connection>
<GID>1386</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1414,619,1414</points>
<connection>
<GID>1527</GID>
<name>OUT_15</name></connection>
<connection>
<GID>1385</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1484</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1404,619,1404</points>
<connection>
<GID>1527</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1390</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1402,619,1402</points>
<connection>
<GID>1527</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>610.5,1392,619,1392</points>
<intersection>610.5 3</intersection>
<intersection>619 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>619,1392,619,1400</points>
<connection>
<GID>1392</GID>
<name>IN_0</name></connection>
<intersection>1392 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>610.5,1392,610.5,1400</points>
<connection>
<GID>1527</GID>
<name>OUT_1</name></connection>
<intersection>1392 1</intersection></vsegment></shape></wire>
<wire>
<ID>1487</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>599,1416,599,1417.5</points>
<connection>
<GID>1526</GID>
<name>count_enable</name></connection>
<connection>
<GID>1402</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>599,1421.5,599,1422.5</points>
<connection>
<GID>1402</GID>
<name>IN_0</name></connection>
<intersection>1422.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>589,1422.5,599,1422.5</points>
<connection>
<GID>1401</GID>
<name>IN_0</name></connection>
<intersection>598 4</intersection>
<intersection>599 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>598,1416,598,1422.5</points>
<connection>
<GID>1526</GID>
<name>load</name></connection>
<intersection>1422.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1489</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600,1416,600,1421.5</points>
<connection>
<GID>1526</GID>
<name>count_up</name></connection>
<connection>
<GID>1403</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1490</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>602,1416,602,1421.5</points>
<connection>
<GID>1526</GID>
<name>carry_out</name></connection>
<connection>
<GID>1404</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1491</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>649.5,1438,649.5,1440.5</points>
<connection>
<GID>1564</GID>
<name>load</name></connection>
<connection>
<GID>1405</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1492</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>667,1480.5,667,1481.5</points>
<connection>
<GID>1458</GID>
<name>load</name></connection>
<connection>
<GID>1406</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1493</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>594.5,1459,594.5,1462.5</points>
<connection>
<GID>1261</GID>
<name>load</name></connection>
<connection>
<GID>1407</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>1494</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1468.5,726,1468.5</points>
<connection>
<GID>1417</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1495</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1470.5,726,1470.5</points>
<connection>
<GID>1416</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1472.5,726,1472.5</points>
<connection>
<GID>1415</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1474.5,726,1474.5</points>
<connection>
<GID>1414</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1498</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1476.5,726,1476.5</points>
<connection>
<GID>1413</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1499</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1478.5,726,1478.5</points>
<connection>
<GID>1412</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1464.5,726,1464.5</points>
<connection>
<GID>1481</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>724.5,1466.5,726,1466.5</points>
<connection>
<GID>1479</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1467.5,726,1467.5</points>
<connection>
<GID>1411</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1469.5,726,1469.5</points>
<connection>
<GID>1410</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1471.5,726,1471.5</points>
<connection>
<GID>1409</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1475.5,726,1475.5</points>
<connection>
<GID>1487</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1477.5,726,1477.5</points>
<connection>
<GID>1486</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1463.5,726,1463.5</points>
<connection>
<GID>1485</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1508</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1465.5,726,1465.5</points>
<connection>
<GID>1483</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1509</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716,1473.5,726,1473.5</points>
<connection>
<GID>1408</GID>
<name>IN_0</name></connection>
<connection>
<GID>1463</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1510</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>745.5,1475.5,748,1475.5</points>
<connection>
<GID>1464</GID>
<name>OUT_12</name></connection>
<connection>
<GID>1427</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1478.5,663,1478.5</points>
<connection>
<GID>1469</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1512</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1476.5,663,1476.5</points>
<connection>
<GID>1471</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1474.5,663,1474.5</points>
<connection>
<GID>1472</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>1514</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1472.5,663,1472.5</points>
<connection>
<GID>1474</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1515</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1470.5,663,1470.5</points>
<connection>
<GID>1475</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1516</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1468.5,663,1468.5</points>
<connection>
<GID>1476</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1466.5,663,1466.5</points>
<connection>
<GID>1431</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1518</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662,1464.5,663,1464.5</points>
<connection>
<GID>1432</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1465.5,663,1465.5</points>
<connection>
<GID>1433</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1463.5,663,1463.5</points>
<connection>
<GID>1434</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1521</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1477.5,663,1477.5</points>
<connection>
<GID>1435</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>1522</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1475.5,663,1475.5</points>
<connection>
<GID>1437</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1523</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1473.5,663,1473.5</points>
<connection>
<GID>1438</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>1524</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1471.5,663,1471.5</points>
<connection>
<GID>1439</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1525</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1469.5,663,1469.5</points>
<connection>
<GID>1440</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>655.5,1467.5,663,1467.5</points>
<connection>
<GID>1441</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>1527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1472.5,696.5,1472.5</points>
<connection>
<GID>1445</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_9</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1472.5,673,1491</points>
<intersection>1472.5 1</intersection>
<intersection>1491 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1491,684,1491</points>
<connection>
<GID>1281</GID>
<name>IN_9</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1528</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1478.5,696.5,1478.5</points>
<connection>
<GID>1442</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_15</name></connection>
<intersection>673 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>673,1478.5,673,1497</points>
<intersection>1478.5 1</intersection>
<intersection>1497 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>673,1497,684,1497</points>
<connection>
<GID>1281</GID>
<name>IN_15</name></connection>
<intersection>673 2</intersection></hsegment></shape></wire>
<wire>
<ID>1529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1476.5,696.5,1476.5</points>
<connection>
<GID>1443</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_13</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1476.5,673,1495</points>
<intersection>1476.5 1</intersection>
<intersection>1495 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1495,684,1495</points>
<connection>
<GID>1281</GID>
<name>IN_13</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1530</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1474.5,696.5,1474.5</points>
<connection>
<GID>1444</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_11</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1474.5,673,1493</points>
<intersection>1474.5 1</intersection>
<intersection>1493 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1493,684,1493</points>
<connection>
<GID>1281</GID>
<name>IN_11</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1470.5,696.5,1470.5</points>
<connection>
<GID>1446</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_7</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1470.5,673,1489</points>
<intersection>1470.5 1</intersection>
<intersection>1489 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1489,684,1489</points>
<connection>
<GID>1281</GID>
<name>IN_7</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1532</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1468.5,696.5,1468.5</points>
<connection>
<GID>1447</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_5</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1468.5,673,1487</points>
<intersection>1468.5 1</intersection>
<intersection>1487 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1487,684,1487</points>
<connection>
<GID>1281</GID>
<name>IN_5</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1466.5,696.5,1466.5</points>
<connection>
<GID>1448</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_3</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1466.5,673,1485</points>
<intersection>1466.5 1</intersection>
<intersection>1485 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1485,684,1485</points>
<connection>
<GID>1281</GID>
<name>IN_3</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>673,1464.5,696.5,1464.5</points>
<connection>
<GID>1449</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_1</name></connection>
<intersection>673 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>673,1464.5,673,1483</points>
<intersection>1464.5 1</intersection>
<intersection>1483 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>673,1483,684,1483</points>
<connection>
<GID>1281</GID>
<name>IN_1</name></connection>
<intersection>673 5</intersection></hsegment></shape></wire>
<wire>
<ID>1535</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1477.5,685,1477.5</points>
<connection>
<GID>1450</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_14</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1477.5,673,1496</points>
<intersection>1477.5 0</intersection>
<intersection>1496 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1496,684,1496</points>
<connection>
<GID>1281</GID>
<name>IN_14</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>1536</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1475.5,685,1475.5</points>
<connection>
<GID>1451</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_12</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1475.5,673,1494</points>
<intersection>1475.5 0</intersection>
<intersection>1494 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1494,684,1494</points>
<connection>
<GID>1281</GID>
<name>IN_12</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire>
<wire>
<ID>1537</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>673,1473.5,685,1473.5</points>
<connection>
<GID>1452</GID>
<name>IN_0</name></connection>
<connection>
<GID>1458</GID>
<name>OUT_10</name></connection>
<intersection>673 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>673,1473.5,673,1492</points>
<intersection>1473.5 0</intersection>
<intersection>1492 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>673,1492,684,1492</points>
<connection>
<GID>1281</GID>
<name>IN_10</name></connection>
<intersection>673 4</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>98.6906,2814.85,1652.69,1799.85</PageViewport>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>340,1294</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>340,1297</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>346,1285.5</position>
<gparam>LABEL_TEXT Skocz gdy 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>341.5,1312.5</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>231.5,1328.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC0</lparam></gate>
<gate>
<ID>226</ID>
<type>DE_TO</type>
<position>360.5,1277</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW3</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_SMALL_INVERTER</type>
<position>346.5,1275.5</position>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>340,1281.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>340,1275.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>340,1278.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>231</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>309.5,1326.5</position>
<output>
<ID>A_equal_B</ID>182 </output>
<output>
<ID>A_greater_B</ID>181 </output>
<output>
<ID>A_less_B</ID>183 </output>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_B_0</ID>200 </input>
<input>
<ID>IN_B_1</ID>201 </input>
<input>
<ID>IN_B_2</ID>202 </input>
<input>
<ID>IN_B_3</ID>203 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>232</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>309.5,1309.5</position>
<output>
<ID>A_equal_B</ID>185 </output>
<output>
<ID>A_greater_B</ID>184 </output>
<output>
<ID>A_less_B</ID>188 </output>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_B_0</ID>204 </input>
<input>
<ID>IN_B_1</ID>205 </input>
<input>
<ID>IN_B_2</ID>206 </input>
<input>
<ID>IN_B_3</ID>207 </input>
<input>
<ID>in_A_equal_B</ID>182 </input>
<input>
<ID>in_A_greater_B</ID>181 </input>
<input>
<ID>in_A_less_B</ID>183 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>233</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>309.5,1292.5</position>
<output>
<ID>A_equal_B</ID>214 </output>
<output>
<ID>A_greater_B</ID>237 </output>
<output>
<ID>A_less_B</ID>213 </output>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_B_0</ID>208 </input>
<input>
<ID>IN_B_1</ID>209 </input>
<input>
<ID>IN_B_2</ID>210 </input>
<input>
<ID>IN_B_3</ID>211 </input>
<input>
<ID>in_A_equal_B</ID>185 </input>
<input>
<ID>in_A_greater_B</ID>184 </input>
<input>
<ID>in_A_less_B</ID>188 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>301,1331.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC0</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>301,1329.5</position>
<input>
<ID>IN_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC1</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>301,1327.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC2</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>301,1325.5</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC3</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>231.5,1326</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC1</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>301,1314.5</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC4</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>231.5,1324</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC2</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>301,1312.5</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC5</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>301,1310.5</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC6</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>301,1308.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC7</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>301,1297.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC8</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>301,1295.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC9</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>301,1293.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC10</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>301,1291.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC11</lparam></gate>
<gate>
<ID>248</ID>
<type>DE_TO</type>
<position>323,1263</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok></lparam></gate>
<gate>
<ID>249</ID>
<type>DE_TO</type>
<position>323,1259</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok=</lparam></gate>
<gate>
<ID>252</ID>
<type>DE_TO</type>
<position>323,1255</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_SMALL_INVERTER</type>
<position>346.5,1316</position>
<input>
<ID>IN_0</ID>178 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_SMALL_INVERTER</type>
<position>346.5,1319.5</position>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>341.5,1322.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>341.5,1316</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B10</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>341.5,1319.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B11</lparam></gate>
<gate>
<ID>258</ID>
<type>DA_FROM</type>
<position>253,1312.5</position>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID COMP0/AddSub1</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_SMALL_INVERTER</type>
<position>256,1276.5</position>
<input>
<ID>IN_0</ID>368 </input>
<output>
<ID>OUT_0</ID>369 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>260</ID>
<type>DE_TO</type>
<position>276.5,1299</position>
<input>
<ID>IN_0</ID>827 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>261</ID>
<type>DE_TO</type>
<position>270,1298</position>
<input>
<ID>IN_0</ID>828 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>186.5,1295</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR6</lparam></gate>
<gate>
<ID>263</ID>
<type>DE_TO</type>
<position>276.5,1297</position>
<input>
<ID>IN_0</ID>826 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>264</ID>
<type>DA_FROM</type>
<position>186.5,1293</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR7</lparam></gate>
<gate>
<ID>265</ID>
<type>DE_TO</type>
<position>270,1296</position>
<input>
<ID>IN_0</ID>824 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>266</ID>
<type>DA_FROM</type>
<position>186.5,1281</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR8</lparam></gate>
<gate>
<ID>267</ID>
<type>DE_TO</type>
<position>276.5,1295</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A4</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>186.5,1279</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR9</lparam></gate>
<gate>
<ID>270</ID>
<type>DE_TO</type>
<position>270,1294</position>
<input>
<ID>IN_0</ID>829 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A5</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>186.5,1277</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR10</lparam></gate>
<gate>
<ID>272</ID>
<type>DE_TO</type>
<position>276.5,1293</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A6</lparam></gate>
<gate>
<ID>668</ID>
<type>DA_FROM</type>
<position>186.5,1258.5</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR14</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>231.5,1267.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC15</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>186.5,1275</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR11</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>186.5,1256.5</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR15</lparam></gate>
<gate>
<ID>286</ID>
<type>DE_TO</type>
<position>270,1292</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A7</lparam></gate>
<gate>
<ID>287</ID>
<type>DE_TO</type>
<position>276.5,1291</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A8</lparam></gate>
<gate>
<ID>288</ID>
<type>DE_TO</type>
<position>270,1290</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A9</lparam></gate>
<gate>
<ID>289</ID>
<type>DE_TO</type>
<position>276.5,1289</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A10</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>231.5,1321.5</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC3</lparam></gate>
<gate>
<ID>291</ID>
<type>DE_TO</type>
<position>270,1288</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A11</lparam></gate>
<gate>
<ID>292</ID>
<type>DE_TO</type>
<position>276.5,1287</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A12</lparam></gate>
<gate>
<ID>293</ID>
<type>DA_FROM</type>
<position>231.5,1310.5</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC4</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>186.5,1262.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR12</lparam></gate>
<gate>
<ID>295</ID>
<type>DE_TO</type>
<position>270,1286</position>
<input>
<ID>IN_0</ID>690 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A13</lparam></gate>
<gate>
<ID>296</ID>
<type>DE_TO</type>
<position>276.5,1285</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A14</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>231.5,1270</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC14</lparam></gate>
<gate>
<ID>299</ID>
<type>DA_FROM</type>
<position>186.5,1260.5</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR13</lparam></gate>
<gate>
<ID>300</ID>
<type>DE_TO</type>
<position>270,1284</position>
<input>
<ID>IN_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A15</lparam></gate>
<gate>
<ID>691</ID>
<type>DA_FROM</type>
<position>231.5,1306</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC6</lparam></gate>
<gate>
<ID>692</ID>
<type>AI_XOR2</type>
<position>220,1324</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>693</ID>
<type>AI_XOR2</type>
<position>220,1319.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>DA_FROM</type>
<position>231.5,1303.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC7</lparam></gate>
<gate>
<ID>696</ID>
<type>AI_XOR2</type>
<position>220,1315</position>
<input>
<ID>IN_0</ID>265 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>697</ID>
<type>AI_XOR2</type>
<position>220,1310.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>698</ID>
<type>AI_XOR2</type>
<position>220,1305.5</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>700</ID>
<type>AI_XOR2</type>
<position>220,1301</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>701</ID>
<type>AI_XOR2</type>
<position>220,1296.5</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>702</ID>
<type>HA_JUNC_2</type>
<position>256,1307</position>
<input>
<ID>N_in0</ID>368 </input>
<input>
<ID>N_in1</ID>367 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>703</ID>
<type>AI_XOR2</type>
<position>220,1292</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>704</ID>
<type>AI_XOR2</type>
<position>220,1287.5</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>705</ID>
<type>AI_XOR2</type>
<position>220,1283</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>706</ID>
<type>AI_XOR2</type>
<position>220,1278.5</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>707</ID>
<type>DA_FROM</type>
<position>232,1292.5</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC8</lparam></gate>
<gate>
<ID>708</ID>
<type>AI_XOR2</type>
<position>220,1274</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>232,1290</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC9</lparam></gate>
<gate>
<ID>710</ID>
<type>AI_XOR2</type>
<position>220,1265</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>DA_FROM</type>
<position>231.5,1308</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC5</lparam></gate>
<gate>
<ID>711</ID>
<type>DA_FROM</type>
<position>232,1288</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC10</lparam></gate>
<gate>
<ID>712</ID>
<type>AI_XOR2</type>
<position>220,1269.5</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>713</ID>
<type>AI_XOR2</type>
<position>220,1260.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>714</ID>
<type>DA_FROM</type>
<position>232,1285.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC11</lparam></gate>
<gate>
<ID>715</ID>
<type>AI_XOR2</type>
<position>220,1256</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>716</ID>
<type>DA_FROM</type>
<position>186.5,1324</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC0</lparam></gate>
<gate>
<ID>717</ID>
<type>DA_FROM</type>
<position>211,1331.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Subt X</lparam></gate>
<gate>
<ID>718</ID>
<type>DA_FROM</type>
<position>210.5,1325</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR0</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>186.5,1322</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC1</lparam></gate>
<gate>
<ID>720</ID>
<type>DA_FROM</type>
<position>210.5,1320.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR1</lparam></gate>
<gate>
<ID>721</ID>
<type>DA_FROM</type>
<position>186.5,1320</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC2</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,1321.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>199 </input>
<input>
<ID>IN_2</ID>219 </input>
<input>
<ID>IN_3</ID>220 </input>
<input>
<ID>IN_B_0</ID>244 </input>
<input>
<ID>IN_B_1</ID>245 </input>
<input>
<ID>IN_B_2</ID>246 </input>
<input>
<ID>IN_B_3</ID>247 </input>
<output>
<ID>OUT_0</ID>277 </output>
<output>
<ID>OUT_1</ID>278 </output>
<output>
<ID>OUT_2</ID>279 </output>
<output>
<ID>OUT_3</ID>280 </output>
<input>
<ID>carry_in</ID>260 </input>
<output>
<ID>carry_out</ID>165 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>722</ID>
<type>DA_FROM</type>
<position>280,1326</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LoadI</lparam></gate>
<gate>
<ID>723</ID>
<type>DA_FROM</type>
<position>210.5,1316</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR2</lparam></gate>
<gate>
<ID>724</ID>
<type>DA_FROM</type>
<position>186.5,1318</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC3</lparam></gate>
<gate>
<ID>725</ID>
<type>DA_FROM</type>
<position>231.5,1274.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC12</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>278.5,1310</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AddI X</lparam></gate>
<gate>
<ID>726</ID>
<type>DA_FROM</type>
<position>186.5,1307</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC4</lparam></gate>
<gate>
<ID>727</ID>
<type>DA_FROM</type>
<position>210.5,1311.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR3</lparam></gate>
<gate>
<ID>728</ID>
<type>AA_TOGGLE</type>
<position>264,1334.5</position>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>309.5,1275</position>
<output>
<ID>A_equal_B</ID>239 </output>
<output>
<ID>A_less_B</ID>238 </output>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>176 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>176 </input>
<input>
<ID>IN_B_0</ID>240 </input>
<input>
<ID>IN_B_1</ID>241 </input>
<input>
<ID>IN_B_2</ID>242 </input>
<input>
<ID>IN_B_3</ID>243 </input>
<input>
<ID>in_A_equal_B</ID>214 </input>
<input>
<ID>in_A_greater_B</ID>237 </input>
<input>
<ID>in_A_less_B</ID>213 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>729</ID>
<type>DA_FROM</type>
<position>210.5,1306.5</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR4</lparam></gate>
<gate>
<ID>730</ID>
<type>DA_FROM</type>
<position>210.5,1302</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR5</lparam></gate>
<gate>
<ID>731</ID>
<type>DA_FROM</type>
<position>186.5,1305</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC5</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>210.5,1297.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR6</lparam></gate>
<gate>
<ID>733</ID>
<type>AI_XOR2</type>
<position>315.5,1263</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,1303.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>222 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>224 </input>
<input>
<ID>IN_B_0</ID>248 </input>
<input>
<ID>IN_B_1</ID>249 </input>
<input>
<ID>IN_B_2</ID>250 </input>
<input>
<ID>IN_B_3</ID>251 </input>
<output>
<ID>OUT_0</ID>281 </output>
<output>
<ID>OUT_1</ID>282 </output>
<output>
<ID>OUT_2</ID>283 </output>
<output>
<ID>OUT_3</ID>284 </output>
<input>
<ID>carry_in</ID>165 </input>
<output>
<ID>carry_out</ID>158 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>736</ID>
<type>DA_FROM</type>
<position>210.5,1293</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR7</lparam></gate>
<gate>
<ID>158</ID>
<type>DE_OR8</type>
<position>265.5,1314</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>216 </input>
<input>
<ID>IN_2</ID>217 </input>
<input>
<ID>IN_3</ID>218 </input>
<input>
<ID>IN_4</ID>260 </input>
<input>
<ID>IN_5</ID>234 </input>
<input>
<ID>IN_6</ID>235 </input>
<input>
<ID>IN_7</ID>236 </input>
<output>
<ID>OUT</ID>367 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>278,1318.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALUS</lparam></gate>
<gate>
<ID>738</ID>
<type>DA_FROM</type>
<position>210.5,1288.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR8</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>279.5,1322</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SkipCond1</lparam></gate>
<gate>
<ID>739</ID>
<type>DA_FROM</type>
<position>301.5,1276.5</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC14</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,1285.5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>227 </input>
<input>
<ID>IN_2</ID>228 </input>
<input>
<ID>IN_3</ID>229 </input>
<input>
<ID>IN_B_0</ID>252 </input>
<input>
<ID>IN_B_1</ID>253 </input>
<input>
<ID>IN_B_2</ID>254 </input>
<input>
<ID>IN_B_3</ID>255 </input>
<output>
<ID>OUT_0</ID>285 </output>
<output>
<ID>OUT_1</ID>286 </output>
<output>
<ID>OUT_2</ID>287 </output>
<output>
<ID>OUT_3</ID>288 </output>
<input>
<ID>carry_in</ID>158 </input>
<output>
<ID>carry_out</ID>159 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>301.5,1274</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC15</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_FULLADDER_4BIT</type>
<position>240,1267.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<input>
<ID>IN_2</ID>232 </input>
<input>
<ID>IN_3</ID>233 </input>
<input>
<ID>IN_B_0</ID>256 </input>
<input>
<ID>IN_B_1</ID>257 </input>
<input>
<ID>IN_B_2</ID>258 </input>
<input>
<ID>IN_B_3</ID>259 </input>
<output>
<ID>OUT_0</ID>289 </output>
<output>
<ID>OUT_1</ID>290 </output>
<output>
<ID>OUT_2</ID>291 </output>
<output>
<ID>OUT_3</ID>292 </output>
<input>
<ID>carry_in</ID>159 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>741</ID>
<type>DA_FROM</type>
<position>301.5,1281</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC12</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>278.5,1313</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Add X</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>301.5,1278.5</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC13</lparam></gate>
<gate>
<ID>164</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>194.5,1264</position>
<output>
<ID>A_equal_B</ID>365 </output>
<output>
<ID>A_greater_B</ID>366 </output>
<output>
<ID>A_less_B</ID>364 </output>
<input>
<ID>IN_0</ID>344 </input>
<input>
<ID>IN_1</ID>345 </input>
<input>
<ID>IN_2</ID>346 </input>
<input>
<ID>IN_3</ID>347 </input>
<input>
<ID>IN_B_0</ID>326 </input>
<input>
<ID>IN_B_1</ID>327 </input>
<input>
<ID>IN_B_2</ID>341 </input>
<input>
<ID>IN_B_3</ID>343 </input>
<input>
<ID>in_A_equal_B</ID>297 </input>
<input>
<ID>in_A_greater_B</ID>296 </input>
<input>
<ID>in_A_less_B</ID>298 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>186.5,1303</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC6</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>278,1315.5</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Load X</lparam></gate>
<gate>
<ID>744</ID>
<type>DA_FROM</type>
<position>210.5,1284</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR9</lparam></gate>
<gate>
<ID>166</ID>
<type>DA_FROM</type>
<position>186.5,1316</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR0</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>210.5,1279.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR10</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>186.5,1314</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR1</lparam></gate>
<gate>
<ID>746</ID>
<type>DA_FROM</type>
<position>210.5,1275</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR11</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND4</type>
<position>354.5,1318.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_2</ID>156 </input>
<input>
<ID>IN_3</ID>160 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>747</ID>
<type>DA_FROM</type>
<position>210.5,1270.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR12</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND4</type>
<position>353,1296</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>161 </input>
<input>
<ID>IN_3</ID>164 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>748</ID>
<type>DA_FROM</type>
<position>186.5,1301</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC7</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>186.5,1312</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR2</lparam></gate>
<gate>
<ID>749</ID>
<type>DA_FROM</type>
<position>186.5,1289</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC8</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>349.5,1327</position>
<gparam>LABEL_TEXT Skocz gdy  0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>750</ID>
<type>DA_FROM</type>
<position>186.5,1287</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC9</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>210.5,1266</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR13</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>186.5,1285</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC10</lparam></gate>
<gate>
<ID>753</ID>
<type>DA_FROM</type>
<position>186.5,1283</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC11</lparam></gate>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>210.5,1261.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR14</lparam></gate>
<gate>
<ID>755</ID>
<type>DA_FROM</type>
<position>210.5,1257</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR15</lparam></gate>
<gate>
<ID>756</ID>
<type>DA_FROM</type>
<position>186.5,1270.5</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC12</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>340,1272.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok></lparam></gate>
<gate>
<ID>757</ID>
<type>DA_FROM</type>
<position>186.5,1268.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC13</lparam></gate>
<gate>
<ID>758</ID>
<type>DA_FROM</type>
<position>231.5,1272</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC13</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>186.5,1310</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR3</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>186.5,1266.5</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC14</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_AND4</type>
<position>354,1277</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>174 </input>
<input>
<ID>IN_3</ID>173 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>760</ID>
<type>DA_FROM</type>
<position>186.5,1264.5</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC15</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>361.5,1318.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW1</lparam></gate>
<gate>
<ID>761</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>264,1291.5</position>
<input>
<ID>ENABLE_0</ID>367 </input>
<input>
<ID>IN_0</ID>363 </input>
<input>
<ID>IN_1</ID>362 </input>
<input>
<ID>IN_10</ID>353 </input>
<input>
<ID>IN_11</ID>352 </input>
<input>
<ID>IN_12</ID>351 </input>
<input>
<ID>IN_13</ID>350 </input>
<input>
<ID>IN_14</ID>349 </input>
<input>
<ID>IN_15</ID>348 </input>
<input>
<ID>IN_2</ID>360 </input>
<input>
<ID>IN_3</ID>361 </input>
<input>
<ID>IN_4</ID>359 </input>
<input>
<ID>IN_5</ID>357 </input>
<input>
<ID>IN_6</ID>358 </input>
<input>
<ID>IN_7</ID>356 </input>
<input>
<ID>IN_8</ID>355 </input>
<input>
<ID>IN_9</ID>354 </input>
<output>
<ID>OUT_0</ID>823 </output>
<output>
<ID>OUT_1</ID>748 </output>
<output>
<ID>OUT_10</ID>829 </output>
<output>
<ID>OUT_11</ID>825 </output>
<output>
<ID>OUT_12</ID>824 </output>
<output>
<ID>OUT_13</ID>826 </output>
<output>
<ID>OUT_14</ID>828 </output>
<output>
<ID>OUT_15</ID>827 </output>
<output>
<ID>OUT_2</ID>690 </output>
<output>
<ID>OUT_3</ID>541 </output>
<output>
<ID>OUT_4</ID>539 </output>
<output>
<ID>OUT_5</ID>374 </output>
<output>
<ID>OUT_6</ID>373 </output>
<output>
<ID>OUT_7</ID>372 </output>
<output>
<ID>OUT_8</ID>371 </output>
<output>
<ID>OUT_9</ID>370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>183</ID>
<type>DA_FROM</type>
<position>186.5,1299</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR4</lparam></gate>
<gate>
<ID>762</ID>
<type>BI_TRI_STATE_4BIT</type>
<position>256,1267.5</position>
<input>
<ID>ENABLE_0</ID>369 </input>
<input>
<ID>IN_0</ID>364 </input>
<input>
<ID>IN_1</ID>365 </input>
<input>
<ID>IN_2</ID>366 </input>
<output>
<ID>OUT_0</ID>348 </output>
<output>
<ID>OUT_1</ID>349 </output>
<output>
<ID>OUT_2</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>346,1304</position>
<gparam>LABEL_TEXT Skocz gdy 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>763</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>256,1291.5</position>
<input>
<ID>ENABLE_0</ID>368 </input>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>291 </input>
<input>
<ID>IN_10</ID>282 </input>
<input>
<ID>IN_11</ID>281 </input>
<input>
<ID>IN_12</ID>280 </input>
<input>
<ID>IN_13</ID>279 </input>
<input>
<ID>IN_14</ID>278 </input>
<input>
<ID>IN_15</ID>277 </input>
<input>
<ID>IN_2</ID>290 </input>
<input>
<ID>IN_3</ID>289 </input>
<input>
<ID>IN_4</ID>288 </input>
<input>
<ID>IN_5</ID>287 </input>
<input>
<ID>IN_6</ID>286 </input>
<input>
<ID>IN_7</ID>285 </input>
<input>
<ID>IN_8</ID>284 </input>
<input>
<ID>IN_9</ID>283 </input>
<output>
<ID>OUT_0</ID>363 </output>
<output>
<ID>OUT_1</ID>362 </output>
<output>
<ID>OUT_10</ID>353 </output>
<output>
<ID>OUT_11</ID>352 </output>
<output>
<ID>OUT_12</ID>351 </output>
<output>
<ID>OUT_13</ID>350 </output>
<output>
<ID>OUT_14</ID>349 </output>
<output>
<ID>OUT_15</ID>348 </output>
<output>
<ID>OUT_2</ID>360 </output>
<output>
<ID>OUT_3</ID>361 </output>
<output>
<ID>OUT_4</ID>359 </output>
<output>
<ID>OUT_5</ID>357 </output>
<output>
<ID>OUT_6</ID>358 </output>
<output>
<ID>OUT_7</ID>356 </output>
<output>
<ID>OUT_8</ID>355 </output>
<output>
<ID>OUT_9</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>185</ID>
<type>FF_GND</type>
<position>295.5,1265</position>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>764</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>194.5,1317.5</position>
<output>
<ID>A_equal_B</ID>300 </output>
<output>
<ID>A_greater_B</ID>299 </output>
<output>
<ID>A_less_B</ID>301 </output>
<input>
<ID>IN_0</ID>306 </input>
<input>
<ID>IN_1</ID>307 </input>
<input>
<ID>IN_2</ID>308 </input>
<input>
<ID>IN_3</ID>309 </input>
<input>
<ID>IN_B_0</ID>302 </input>
<input>
<ID>IN_B_1</ID>303 </input>
<input>
<ID>IN_B_2</ID>304 </input>
<input>
<ID>IN_B_3</ID>305 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>186</ID>
<type>DA_FROM</type>
<position>186.5,1297</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MDR5</lparam></gate>
<gate>
<ID>765</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>194.5,1300</position>
<output>
<ID>A_equal_B</ID>294 </output>
<output>
<ID>A_greater_B</ID>293 </output>
<output>
<ID>A_less_B</ID>295 </output>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>315 </input>
<input>
<ID>IN_2</ID>316 </input>
<input>
<ID>IN_3</ID>317 </input>
<input>
<ID>IN_B_0</ID>310 </input>
<input>
<ID>IN_B_1</ID>311 </input>
<input>
<ID>IN_B_2</ID>312 </input>
<input>
<ID>IN_B_3</ID>313 </input>
<input>
<ID>in_A_equal_B</ID>300 </input>
<input>
<ID>in_A_greater_B</ID>299 </input>
<input>
<ID>in_A_less_B</ID>301 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>187</ID>
<type>DA_FROM</type>
<position>340,1291</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Skok=</lparam></gate>
<gate>
<ID>766</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>194.5,1282</position>
<output>
<ID>A_equal_B</ID>297 </output>
<output>
<ID>A_greater_B</ID>296 </output>
<output>
<ID>A_less_B</ID>298 </output>
<input>
<ID>IN_0</ID>322 </input>
<input>
<ID>IN_1</ID>323 </input>
<input>
<ID>IN_2</ID>324 </input>
<input>
<ID>IN_3</ID>325 </input>
<input>
<ID>IN_B_0</ID>318 </input>
<input>
<ID>IN_B_1</ID>319 </input>
<input>
<ID>IN_B_2</ID>320 </input>
<input>
<ID>IN_B_3</ID>321 </input>
<input>
<ID>in_A_equal_B</ID>294 </input>
<input>
<ID>in_A_greater_B</ID>293 </input>
<input>
<ID>in_A_less_B</ID>295 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>359.5,1296</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PCW2</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_SMALL_INVERTER</type>
<position>345,1297</position>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>340,1300</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SkipCond</lparam></gate>
<wire>
<ID>823</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1284,268,1284</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1296,268,1296</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1295,274.5,1295</points>
<connection>
<GID>761</GID>
<name>OUT_11</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1297,274.5,1297</points>
<connection>
<GID>761</GID>
<name>OUT_13</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1299,274.5,1299</points>
<connection>
<GID>761</GID>
<name>OUT_15</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1298,268,1298</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1294,268,1294</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>539</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1288,268,1288</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1287,274.5,1287</points>
<connection>
<GID>761</GID>
<name>OUT_3</name></connection>
<connection>
<GID>292</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,1322.5,351.5,1322.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>351.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>351.5,1321.5,351.5,1322.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>1322.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>348.5,1319.5,351.5,1319.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<connection>
<GID>168</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,1316,350,1317.5</points>
<intersection>1316 2</intersection>
<intersection>1317.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,1317.5,351.5,1317.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,1316,350,1316</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>357.5,1318.5,359.5,1318.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,1293.5,239,1295.5</points>
<connection>
<GID>161</GID>
<name>carry_in</name></connection>
<connection>
<GID>157</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,1275.5,239,1277.5</points>
<connection>
<GID>162</GID>
<name>carry_in</name></connection>
<connection>
<GID>161</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>351,1312.5,351,1315.5</points>
<intersection>1312.5 2</intersection>
<intersection>1315.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>351,1315.5,351.5,1315.5</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>351 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>343.5,1312.5,351,1312.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>351 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,1294,350,1295</points>
<connection>
<GID>169</GID>
<name>IN_2</name></connection>
<intersection>1294 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>342,1294,350,1294</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>347,1297,350,1297</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>342,1300,350,1300</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>350 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>350,1299,350,1300</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>1300 1</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,1291,349.5,1293</points>
<intersection>1291 2</intersection>
<intersection>1293 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>349.5,1293,350,1293</points>
<connection>
<GID>169</GID>
<name>IN_3</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,1291,349.5,1291</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>239,1311.5,239,1313.5</points>
<connection>
<GID>157</GID>
<name>carry_in</name></connection>
<connection>
<GID>143</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1319.5,225,1324</points>
<intersection>1319.5 1</intersection>
<intersection>1324 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1319.5,236,1319.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1324,225,1324</points>
<connection>
<GID>692</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>356,1296,357.5,1296</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>349.5,1280,349.5,1281.5</points>
<intersection>1280 3</intersection>
<intersection>1281.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>342,1281.5,349.5,1281.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>349.5,1280,351,1280</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>349.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>357,1277,358.5,1277</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,1272.5,350,1274</points>
<intersection>1272.5 2</intersection>
<intersection>1274 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,1274,351,1274</points>
<connection>
<GID>181</GID>
<name>IN_3</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,1272.5,350,1272.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,1275.5,350,1276</points>
<intersection>1275.5 2</intersection>
<intersection>1276 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,1276,351,1276</points>
<connection>
<GID>181</GID>
<name>IN_2</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>348.5,1275.5,350,1275.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,1278,350,1278.5</points>
<intersection>1278 1</intersection>
<intersection>1278.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,1278,351,1278</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,1278.5,350,1278.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295.5,1266,295.5,1324.5</points>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection>
<intersection>1270 33</intersection>
<intersection>1271 34</intersection>
<intersection>1272 35</intersection>
<intersection>1273 26</intersection>
<intersection>1287.5 27</intersection>
<intersection>1288.5 28</intersection>
<intersection>1289.5 29</intersection>
<intersection>1290.5 14</intersection>
<intersection>1304.5 15</intersection>
<intersection>1305.5 16</intersection>
<intersection>1306.5 17</intersection>
<intersection>1307.5 6</intersection>
<intersection>1321.5 7</intersection>
<intersection>1322.5 8</intersection>
<intersection>1323.5 9</intersection>
<intersection>1324.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295.5,1324.5,305.5,1324.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>295.5,1307.5,305.5,1307.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>295.5,1321.5,305.5,1321.5</points>
<connection>
<GID>231</GID>
<name>IN_3</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>295.5,1322.5,305.5,1322.5</points>
<connection>
<GID>231</GID>
<name>IN_2</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>295.5,1323.5,305.5,1323.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>295.5,1290.5,305.5,1290.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>295.5,1304.5,305.5,1304.5</points>
<connection>
<GID>232</GID>
<name>IN_3</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>295.5,1305.5,305.5,1305.5</points>
<connection>
<GID>232</GID>
<name>IN_2</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>295.5,1306.5,305.5,1306.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>295.5,1273,305.5,1273</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>295.5,1287.5,305.5,1287.5</points>
<connection>
<GID>233</GID>
<name>IN_3</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>295.5,1288.5,305.5,1288.5</points>
<connection>
<GID>233</GID>
<name>IN_2</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>295.5,1289.5,305.5,1289.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>295.5,1270,305.5,1270</points>
<connection>
<GID>150</GID>
<name>IN_3</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>295.5,1271,305.5,1271</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>295.5 0</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>295.5,1272,305.5,1272</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>295.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,1319.5,344.5,1319.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>257</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343.5,1316,344.5,1316</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>256</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>342,1297,343,1297</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>191</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>342,1275.5,344.5,1275.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,1317.5,307.5,1318.5</points>
<connection>
<GID>232</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>231</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,1317.5,309.5,1318.5</points>
<connection>
<GID>232</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>231</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,1317.5,311.5,1318.5</points>
<connection>
<GID>232</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>231</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,1300.5,307.5,1301.5</points>
<connection>
<GID>233</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>232</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,1300.5,309.5,1301.5</points>
<connection>
<GID>233</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>232</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,1300.5,311.5,1301.5</points>
<connection>
<GID>233</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>232</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,1318.5,224,1319.5</points>
<intersection>1318.5 1</intersection>
<intersection>1319.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,1318.5,236,1318.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1319.5,224,1319.5</points>
<connection>
<GID>693</GID>
<name>OUT</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>303,1331.5,305.5,1331.5</points>
<connection>
<GID>231</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1329.5,304.5,1330.5</points>
<intersection>1329.5 2</intersection>
<intersection>1330.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1330.5,305.5,1330.5</points>
<connection>
<GID>231</GID>
<name>IN_B_1</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1329.5,304.5,1329.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1327.5,304.5,1329.5</points>
<intersection>1327.5 2</intersection>
<intersection>1329.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1329.5,305.5,1329.5</points>
<connection>
<GID>231</GID>
<name>IN_B_2</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1327.5,304.5,1327.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1325.5,304.5,1328.5</points>
<intersection>1325.5 2</intersection>
<intersection>1328.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1328.5,305.5,1328.5</points>
<connection>
<GID>231</GID>
<name>IN_B_3</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1325.5,304.5,1325.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>303,1314.5,305.5,1314.5</points>
<connection>
<GID>232</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>303,1313.5,305.5,1313.5</points>
<connection>
<GID>232</GID>
<name>IN_B_1</name></connection>
<intersection>303 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>303,1312.5,303,1313.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>1313.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1310.5,304.5,1312.5</points>
<intersection>1310.5 2</intersection>
<intersection>1312.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1312.5,305.5,1312.5</points>
<connection>
<GID>232</GID>
<name>IN_B_2</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1310.5,304.5,1310.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1308.5,304.5,1311.5</points>
<intersection>1308.5 2</intersection>
<intersection>1311.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1311.5,305.5,1311.5</points>
<connection>
<GID>232</GID>
<name>IN_B_3</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1308.5,304.5,1308.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>303,1297.5,305.5,1297.5</points>
<connection>
<GID>233</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1295.5,304.5,1296.5</points>
<intersection>1295.5 2</intersection>
<intersection>1296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1296.5,305.5,1296.5</points>
<connection>
<GID>233</GID>
<name>IN_B_1</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1295.5,304.5,1295.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1293.5,304.5,1295.5</points>
<intersection>1293.5 2</intersection>
<intersection>1295.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1295.5,305.5,1295.5</points>
<connection>
<GID>233</GID>
<name>IN_B_2</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1293.5,304.5,1293.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1291.5,304.5,1294.5</points>
<intersection>1291.5 2</intersection>
<intersection>1294.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304.5,1294.5,305.5,1294.5</points>
<connection>
<GID>233</GID>
<name>IN_B_3</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>303,1291.5,304.5,1291.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>318.5,1263,321,1263</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<connection>
<GID>733</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,1283,311.5,1284.5</points>
<connection>
<GID>150</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>233</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,1283,309.5,1284.5</points>
<connection>
<GID>150</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>233</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,1310,273.5,1310.5</points>
<intersection>1310 2</intersection>
<intersection>1310.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1310.5,273.5,1310.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>273.5,1310,276.5,1310</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>273.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273.5,1311.5,273.5,1313</points>
<intersection>1311.5 1</intersection>
<intersection>1313 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1311.5,273.5,1311.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>273.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>273.5,1313,276.5,1313</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>273.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,1312.5,273,1315.5</points>
<intersection>1312.5 1</intersection>
<intersection>1315.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1312.5,273,1312.5</points>
<connection>
<GID>158</GID>
<name>IN_2</name></connection>
<intersection>273 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>273,1315.5,276,1315.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,1313.5,272.5,1318.5</points>
<intersection>1313.5 1</intersection>
<intersection>1318.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1313.5,272.5,1313.5</points>
<connection>
<GID>158</GID>
<name>IN_3</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>272.5,1318.5,276,1318.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,1315,224,1317.5</points>
<intersection>1315 2</intersection>
<intersection>1317.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,1317.5,236,1317.5</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1315,224,1315</points>
<connection>
<GID>696</GID>
<name>OUT</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1310.5,225,1316.5</points>
<intersection>1310.5 2</intersection>
<intersection>1316.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1316.5,236,1316.5</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1310.5,225,1310.5</points>
<connection>
<GID>697</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,1301.5,226,1305.5</points>
<intersection>1301.5 1</intersection>
<intersection>1305.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,1301.5,236,1301.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1305.5,226,1305.5</points>
<connection>
<GID>698</GID>
<name>OUT</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>225,1300.5,236,1300.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>225 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>225,1300.5,225,1301</points>
<intersection>1300.5 1</intersection>
<intersection>1301 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>223,1301,225,1301</points>
<connection>
<GID>700</GID>
<name>OUT</name></connection>
<intersection>225 3</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1296.5,225,1299.5</points>
<intersection>1296.5 2</intersection>
<intersection>1299.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1299.5,236,1299.5</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1296.5,225,1296.5</points>
<connection>
<GID>701</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>226,1292,226,1298.5</points>
<intersection>1292 2</intersection>
<intersection>1298.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>226,1298.5,236,1298.5</points>
<connection>
<GID>157</GID>
<name>IN_3</name></connection>
<intersection>226 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1292,226,1292</points>
<connection>
<GID>703</GID>
<name>OUT</name></connection>
<intersection>226 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1283.5,225,1287.5</points>
<intersection>1283.5 1</intersection>
<intersection>1287.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1283.5,236,1283.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1287.5,225,1287.5</points>
<connection>
<GID>704</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>224,1282.5,236,1282.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>224 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>224,1282.5,224,1283</points>
<intersection>1282.5 1</intersection>
<intersection>1283 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>223,1283,224,1283</points>
<connection>
<GID>705</GID>
<name>OUT</name></connection>
<intersection>224 3</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,1278.5,224,1281.5</points>
<intersection>1278.5 2</intersection>
<intersection>1281.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,1281.5,236,1281.5</points>
<connection>
<GID>161</GID>
<name>IN_2</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1278.5,224,1278.5</points>
<connection>
<GID>706</GID>
<name>OUT</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1274,225,1280.5</points>
<intersection>1274 2</intersection>
<intersection>1280.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1280.5,236,1280.5</points>
<connection>
<GID>161</GID>
<name>IN_3</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1274,225,1274</points>
<connection>
<GID>708</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1265.5,225,1269.5</points>
<intersection>1265.5 1</intersection>
<intersection>1269.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1265.5,236,1265.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1269.5,225,1269.5</points>
<connection>
<GID>712</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>224,1264.5,236,1264.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>224 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>224,1264.5,224,1265</points>
<intersection>1264.5 1</intersection>
<intersection>1265 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>223,1265,224,1265</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<intersection>224 3</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,1260.5,224,1263.5</points>
<intersection>1260.5 2</intersection>
<intersection>1263.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,1263.5,236,1263.5</points>
<connection>
<GID>162</GID>
<name>IN_2</name></connection>
<intersection>224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1260.5,224,1260.5</points>
<connection>
<GID>713</GID>
<name>OUT</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,1256,225,1262.5</points>
<intersection>1256 2</intersection>
<intersection>1262.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,1262.5,236,1262.5</points>
<connection>
<GID>162</GID>
<name>IN_3</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,1256,225,1256</points>
<connection>
<GID>715</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270,1316.5,270,1334.5</points>
<intersection>1316.5 1</intersection>
<intersection>1334.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1316.5,270,1316.5</points>
<connection>
<GID>158</GID>
<name>IN_5</name></connection>
<intersection>270 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266,1334.5,270,1334.5</points>
<connection>
<GID>728</GID>
<name>OUT_0</name></connection>
<intersection>270 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>271,1315.5,271,1326</points>
<intersection>1315.5 1</intersection>
<intersection>1326 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268.5,1315.5,271,1315.5</points>
<connection>
<GID>158</GID>
<name>IN_6</name></connection>
<intersection>271 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>271,1326,278,1326</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<intersection>271 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272,1314.5,272,1322</points>
<intersection>1314.5 2</intersection>
<intersection>1322 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>272,1322,277.5,1322</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>272 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>268.5,1314.5,272,1314.5</points>
<connection>
<GID>158</GID>
<name>IN_7</name></connection>
<intersection>272 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>307.5,1283,307.5,1284.5</points>
<connection>
<GID>150</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>233</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>311.5,1264,311.5,1267</points>
<connection>
<GID>150</GID>
<name>A_less_B</name></connection>
<intersection>1264 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>311.5,1264,312.5,1264</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<intersection>311.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309.5,1259,309.5,1267</points>
<connection>
<GID>150</GID>
<name>A_equal_B</name></connection>
<intersection>1259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>309.5,1259,321,1259</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>309.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1280,304.5,1281</points>
<intersection>1280 2</intersection>
<intersection>1281 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,1281,304.5,1281</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,1280,305.5,1280</points>
<connection>
<GID>150</GID>
<name>IN_B_0</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1278.5,304.5,1279</points>
<intersection>1278.5 1</intersection>
<intersection>1279 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,1278.5,304.5,1278.5</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,1279,305.5,1279</points>
<connection>
<GID>150</GID>
<name>IN_B_1</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,1276.5,304,1278</points>
<intersection>1276.5 1</intersection>
<intersection>1278 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,1276.5,304,1276.5</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304,1278,305.5,1278</points>
<connection>
<GID>150</GID>
<name>IN_B_2</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304.5,1255,304.5,1277</points>
<intersection>1255 3</intersection>
<intersection>1262 5</intersection>
<intersection>1274 1</intersection>
<intersection>1277 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>303.5,1274,304.5,1274</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>304.5,1277,305.5,1277</points>
<connection>
<GID>150</GID>
<name>IN_B_3</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>304.5,1255,321,1255</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>304.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>304.5,1262,312.5,1262</points>
<connection>
<GID>733</GID>
<name>IN_1</name></connection>
<intersection>304.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1326.5,235,1328.5</points>
<intersection>1326.5 3</intersection>
<intersection>1328.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1328.5,235,1328.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>235,1326.5,236,1326.5</points>
<connection>
<GID>143</GID>
<name>IN_B_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234,1325.5,236,1325.5</points>
<connection>
<GID>143</GID>
<name>IN_B_1</name></connection>
<intersection>234 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>234,1325.5,234,1326</points>
<intersection>1325.5 1</intersection>
<intersection>1326 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>233.5,1326,234,1326</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>234 6</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>234,1324,234,1324.5</points>
<intersection>1324 6</intersection>
<intersection>1324.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>234,1324.5,236,1324.5</points>
<connection>
<GID>143</GID>
<name>IN_B_2</name></connection>
<intersection>234 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>233.5,1324,234,1324</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>234 4</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>233.5,1321.5,235,1321.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>235 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>235,1321.5,235,1323.5</points>
<intersection>1321.5 2</intersection>
<intersection>1323.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>235,1323.5,236,1323.5</points>
<connection>
<GID>143</GID>
<name>IN_B_3</name></connection>
<intersection>235 4</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1308.5,235,1310.5</points>
<intersection>1308.5 1</intersection>
<intersection>1310.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1308.5,236,1308.5</points>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1310.5,235,1310.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,1307.5,234.5,1308</points>
<intersection>1307.5 1</intersection>
<intersection>1308 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,1307.5,236,1307.5</points>
<connection>
<GID>157</GID>
<name>IN_B_1</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1308,234.5,1308</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,1306,234.5,1306.5</points>
<intersection>1306 2</intersection>
<intersection>1306.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>234.5,1306.5,236,1306.5</points>
<connection>
<GID>157</GID>
<name>IN_B_2</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1306,234.5,1306</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1303.5,235,1305.5</points>
<intersection>1303.5 2</intersection>
<intersection>1305.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1305.5,236,1305.5</points>
<connection>
<GID>157</GID>
<name>IN_B_3</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1303.5,235,1303.5</points>
<connection>
<GID>695</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1290.5,235,1292.5</points>
<intersection>1290.5 1</intersection>
<intersection>1292.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1290.5,236,1290.5</points>
<connection>
<GID>161</GID>
<name>IN_B_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,1292.5,235,1292.5</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1289.5,235,1290</points>
<intersection>1289.5 1</intersection>
<intersection>1290 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1289.5,236,1289.5</points>
<connection>
<GID>161</GID>
<name>IN_B_1</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,1290,235,1290</points>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1288,235,1288.5</points>
<intersection>1288 2</intersection>
<intersection>1288.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1288.5,236,1288.5</points>
<connection>
<GID>161</GID>
<name>IN_B_2</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,1288,235,1288</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1285.5,235,1287.5</points>
<intersection>1285.5 2</intersection>
<intersection>1287.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,1287.5,236,1287.5</points>
<connection>
<GID>161</GID>
<name>IN_B_3</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>234,1285.5,235,1285.5</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1272.5,235,1274.5</points>
<intersection>1272.5 3</intersection>
<intersection>1274.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1274.5,235,1274.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>235,1272.5,236,1272.5</points>
<connection>
<GID>162</GID>
<name>IN_B_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>234,1271.5,236,1271.5</points>
<connection>
<GID>162</GID>
<name>IN_B_1</name></connection>
<intersection>234 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>234,1271.5,234,1272</points>
<intersection>1271.5 2</intersection>
<intersection>1272 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>233.5,1272,234,1272</points>
<connection>
<GID>758</GID>
<name>IN_0</name></connection>
<intersection>234 4</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>234,1270.5,236,1270.5</points>
<connection>
<GID>162</GID>
<name>IN_B_2</name></connection>
<intersection>234 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>234,1270,234,1270.5</points>
<intersection>1270 6</intersection>
<intersection>1270.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>233.5,1270,234,1270</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>234 5</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,1267.5,235,1269.5</points>
<intersection>1267.5 2</intersection>
<intersection>1269.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>233.5,1267.5,235,1267.5</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>235,1269.5,236,1269.5</points>
<connection>
<GID>162</GID>
<name>IN_B_3</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,1255,216,1331.5</points>
<intersection>1255 1</intersection>
<intersection>1259.5 22</intersection>
<intersection>1264 23</intersection>
<intersection>1268.5 24</intersection>
<intersection>1273 21</intersection>
<intersection>1277.5 18</intersection>
<intersection>1282 13</intersection>
<intersection>1286.5 12</intersection>
<intersection>1290.5 11</intersection>
<intersection>1295.5 10</intersection>
<intersection>1300 9</intersection>
<intersection>1304.5 8</intersection>
<intersection>1309.5 7</intersection>
<intersection>1314 6</intersection>
<intersection>1318.5 5</intersection>
<intersection>1323 27</intersection>
<intersection>1331.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>216,1255,217,1255</points>
<connection>
<GID>715</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>213,1331.5,269.5,1331.5</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<intersection>216 0</intersection>
<intersection>239 31</intersection>
<intersection>269.5 29</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>216,1318.5,217,1318.5</points>
<connection>
<GID>693</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>216,1314,217,1314</points>
<connection>
<GID>696</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>216,1309.5,217,1309.5</points>
<connection>
<GID>697</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>216,1304.5,217,1304.5</points>
<connection>
<GID>698</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>216,1300,217,1300</points>
<connection>
<GID>700</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>216,1295.5,217,1295.5</points>
<connection>
<GID>701</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>216,1290.5,217,1290.5</points>
<intersection>216 0</intersection>
<intersection>217 30</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>216,1286.5,217,1286.5</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>216,1282,217,1282</points>
<connection>
<GID>705</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>216,1277.5,217,1277.5</points>
<connection>
<GID>706</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>216,1273,217,1273</points>
<connection>
<GID>708</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>216,1259.5,217,1259.5</points>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>216,1264,217,1264</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>216,1268.5,217,1268.5</points>
<connection>
<GID>712</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>216,1323,217,1323</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<intersection>216 0</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>269.5,1317.5,269.5,1331.5</points>
<intersection>1317.5 32</intersection>
<intersection>1331.5 2</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>217,1290.5,217,1291</points>
<connection>
<GID>703</GID>
<name>IN_1</name></connection>
<intersection>1290.5 11</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>239,1329.5,239,1331.5</points>
<connection>
<GID>143</GID>
<name>carry_in</name></connection>
<intersection>1331.5 2</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>268.5,1317.5,269.5,1317.5</points>
<connection>
<GID>158</GID>
<name>IN_4</name></connection>
<intersection>269.5 29</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1257,217,1257</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<connection>
<GID>715</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1261.5,217,1261.5</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<connection>
<GID>713</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1325,217,1325</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<connection>
<GID>692</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1320.5,217,1320.5</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1316,217,1316</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<connection>
<GID>696</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1311.5,217,1311.5</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1306.5,217,1306.5</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<connection>
<GID>698</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1302,217,1302</points>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<connection>
<GID>700</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1297.5,217,1297.5</points>
<connection>
<GID>732</GID>
<name>IN_0</name></connection>
<connection>
<GID>701</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1293,217,1293</points>
<connection>
<GID>736</GID>
<name>IN_0</name></connection>
<connection>
<GID>703</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1288.5,217,1288.5</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<connection>
<GID>704</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1284,217,1284</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<connection>
<GID>705</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1279.5,217,1279.5</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<connection>
<GID>706</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1275,217,1275</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<connection>
<GID>708</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1270.5,217,1270.5</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<connection>
<GID>712</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>212.5,1266,217,1266</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<connection>
<GID>710</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,1299,251,1323</points>
<intersection>1299 1</intersection>
<intersection>1323 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,1299,254,1299</points>
<connection>
<GID>763</GID>
<name>IN_15</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1323,251,1323</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>251 0</intersection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,1298,250,1322</points>
<intersection>1298 1</intersection>
<intersection>1322 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,1298,254,1298</points>
<connection>
<GID>763</GID>
<name>IN_14</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1322,250,1322</points>
<connection>
<GID>143</GID>
<name>OUT_1</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,1297,249,1321</points>
<intersection>1297 1</intersection>
<intersection>1321 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249,1297,254,1297</points>
<connection>
<GID>763</GID>
<name>IN_13</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1321,249,1321</points>
<connection>
<GID>143</GID>
<name>OUT_2</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,1296,248,1320</points>
<intersection>1296 1</intersection>
<intersection>1320 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,1296,254,1296</points>
<connection>
<GID>763</GID>
<name>IN_12</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1320,248,1320</points>
<connection>
<GID>143</GID>
<name>OUT_3</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,1295,247,1305</points>
<intersection>1295 1</intersection>
<intersection>1305 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,1295,254,1295</points>
<connection>
<GID>763</GID>
<name>IN_11</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1305,247,1305</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,1294,246,1304</points>
<intersection>1294 1</intersection>
<intersection>1304 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246,1294,254,1294</points>
<connection>
<GID>763</GID>
<name>IN_10</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1304,246,1304</points>
<connection>
<GID>157</GID>
<name>OUT_1</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,1293,245,1303</points>
<intersection>1293 1</intersection>
<intersection>1303 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,1293,254,1293</points>
<connection>
<GID>763</GID>
<name>IN_9</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1303,245,1303</points>
<connection>
<GID>157</GID>
<name>OUT_2</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,1292,244,1302</points>
<connection>
<GID>157</GID>
<name>OUT_3</name></connection>
<intersection>1292 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,1292,254,1292</points>
<connection>
<GID>763</GID>
<name>IN_8</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,1287,244,1291</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>1291 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>244,1291,254,1291</points>
<connection>
<GID>763</GID>
<name>IN_7</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245,1286,245,1290</points>
<intersection>1286 2</intersection>
<intersection>1290 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245,1290,254,1290</points>
<connection>
<GID>763</GID>
<name>IN_6</name></connection>
<intersection>245 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1286,245,1286</points>
<connection>
<GID>161</GID>
<name>OUT_1</name></connection>
<intersection>245 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>246,1285,246,1289</points>
<intersection>1285 2</intersection>
<intersection>1289 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>246,1289,254,1289</points>
<connection>
<GID>763</GID>
<name>IN_5</name></connection>
<intersection>246 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1285,246,1285</points>
<connection>
<GID>161</GID>
<name>OUT_2</name></connection>
<intersection>246 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>247,1284,247,1288</points>
<intersection>1284 2</intersection>
<intersection>1288 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>247,1288,254,1288</points>
<connection>
<GID>763</GID>
<name>IN_4</name></connection>
<intersection>247 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1284,247,1284</points>
<connection>
<GID>161</GID>
<name>OUT_3</name></connection>
<intersection>247 0</intersection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>248,1269,248,1287</points>
<intersection>1269 2</intersection>
<intersection>1287 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>248,1287,254,1287</points>
<connection>
<GID>763</GID>
<name>IN_3</name></connection>
<intersection>248 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1269,248,1269</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>248 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249,1268,249,1286</points>
<intersection>1268 2</intersection>
<intersection>1286 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>249,1286,254,1286</points>
<connection>
<GID>763</GID>
<name>IN_2</name></connection>
<intersection>249 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1268,249,1268</points>
<connection>
<GID>162</GID>
<name>OUT_1</name></connection>
<intersection>249 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,1267,250,1285</points>
<intersection>1267 2</intersection>
<intersection>1285 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>250,1285,254,1285</points>
<connection>
<GID>763</GID>
<name>IN_1</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1267,250,1267</points>
<connection>
<GID>162</GID>
<name>OUT_2</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,1266,251,1284</points>
<intersection>1266 2</intersection>
<intersection>1284 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>251,1284,254,1284</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>251 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,1266,251,1266</points>
<connection>
<GID>162</GID>
<name>OUT_3</name></connection>
<intersection>251 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,1290,192.5,1292</points>
<connection>
<GID>766</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>765</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,1290,194.5,1292</points>
<connection>
<GID>766</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>765</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,1290,196.5,1292</points>
<connection>
<GID>766</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>765</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,1272,192.5,1274</points>
<connection>
<GID>164</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>766</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,1272,194.5,1274</points>
<connection>
<GID>164</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>766</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,1272,196.5,1274</points>
<connection>
<GID>164</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>766</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,1308,192.5,1309.5</points>
<connection>
<GID>765</GID>
<name>in_A_greater_B</name></connection>
<connection>
<GID>764</GID>
<name>A_greater_B</name></connection></vsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,1308,194.5,1309.5</points>
<connection>
<GID>765</GID>
<name>in_A_equal_B</name></connection>
<connection>
<GID>764</GID>
<name>A_equal_B</name></connection></vsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,1308,196.5,1309.5</points>
<connection>
<GID>765</GID>
<name>in_A_less_B</name></connection>
<connection>
<GID>764</GID>
<name>A_less_B</name></connection></vsegment></shape></wire>
<wire>
<ID>690</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1286,268,1286</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1322.5,189.5,1324</points>
<intersection>1322.5 1</intersection>
<intersection>1324 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1322.5,190.5,1322.5</points>
<connection>
<GID>764</GID>
<name>IN_B_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1324,189.5,1324</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1321.5,189.5,1322</points>
<intersection>1321.5 1</intersection>
<intersection>1322 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1321.5,190.5,1321.5</points>
<connection>
<GID>764</GID>
<name>IN_B_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1322,189.5,1322</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1320,189.5,1320.5</points>
<intersection>1320 2</intersection>
<intersection>1320.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1320.5,190.5,1320.5</points>
<connection>
<GID>764</GID>
<name>IN_B_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1320,189.5,1320</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1318,189.5,1319.5</points>
<intersection>1318 2</intersection>
<intersection>1319.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1319.5,190.5,1319.5</points>
<connection>
<GID>764</GID>
<name>IN_B_3</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1318,189.5,1318</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1315.5,189.5,1316</points>
<intersection>1315.5 1</intersection>
<intersection>1316 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1315.5,190.5,1315.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1316,189.5,1316</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1314,189.5,1314.5</points>
<intersection>1314 2</intersection>
<intersection>1314.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1314.5,190.5,1314.5</points>
<connection>
<GID>764</GID>
<name>IN_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1314,189.5,1314</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1312,189.5,1313.5</points>
<intersection>1312 2</intersection>
<intersection>1313.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1313.5,190.5,1313.5</points>
<connection>
<GID>764</GID>
<name>IN_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1312,189.5,1312</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1310,190,1312.5</points>
<intersection>1310 2</intersection>
<intersection>1312.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1312.5,190.5,1312.5</points>
<connection>
<GID>764</GID>
<name>IN_3</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1310,190,1310</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1305,190,1307</points>
<intersection>1305 1</intersection>
<intersection>1307 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1305,190.5,1305</points>
<connection>
<GID>765</GID>
<name>IN_B_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1307,190,1307</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1304,189.5,1305</points>
<intersection>1304 1</intersection>
<intersection>1305 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1304,190.5,1304</points>
<connection>
<GID>765</GID>
<name>IN_B_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1305,189.5,1305</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,1303,190.5,1303</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<connection>
<GID>765</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>189,1302,190.5,1302</points>
<connection>
<GID>765</GID>
<name>IN_B_3</name></connection>
<intersection>189 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>189,1301,189,1302</points>
<intersection>1301 10</intersection>
<intersection>1302 6</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>188.5,1301,189,1301</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<intersection>189 9</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1298,189.5,1299</points>
<intersection>1298 1</intersection>
<intersection>1299 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1298,190.5,1298</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1299,189.5,1299</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,1297,190.5,1297</points>
<connection>
<GID>765</GID>
<name>IN_1</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1295,189.5,1296</points>
<intersection>1295 2</intersection>
<intersection>1296 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1296,190.5,1296</points>
<connection>
<GID>765</GID>
<name>IN_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1295,189.5,1295</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1293,190,1295</points>
<intersection>1293 2</intersection>
<intersection>1295 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1295,190.5,1295</points>
<connection>
<GID>765</GID>
<name>IN_3</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1293,190,1293</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1287,190,1289</points>
<intersection>1287 1</intersection>
<intersection>1289 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1287,190.5,1287</points>
<connection>
<GID>766</GID>
<name>IN_B_0</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1289,190,1289</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1286,189.5,1287</points>
<intersection>1286 1</intersection>
<intersection>1287 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1286,190.5,1286</points>
<connection>
<GID>766</GID>
<name>IN_B_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1287,189.5,1287</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,1285,190.5,1285</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<connection>
<GID>766</GID>
<name>IN_B_2</name></connection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1283,189.5,1284</points>
<intersection>1283 2</intersection>
<intersection>1284 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1284,190.5,1284</points>
<connection>
<GID>766</GID>
<name>IN_B_3</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1283,189.5,1283</points>
<connection>
<GID>753</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1280,189.5,1281</points>
<intersection>1280 1</intersection>
<intersection>1281 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1280,190.5,1280</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1281,189.5,1281</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188.5,1279,190.5,1279</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>766</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1277,189.5,1278</points>
<intersection>1277 2</intersection>
<intersection>1278 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1278,190.5,1278</points>
<connection>
<GID>766</GID>
<name>IN_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1277,189.5,1277</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1275,190,1277</points>
<intersection>1275 2</intersection>
<intersection>1277 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1277,190.5,1277</points>
<connection>
<GID>766</GID>
<name>IN_3</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1275,190,1275</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1269,189.5,1270.5</points>
<intersection>1269 1</intersection>
<intersection>1270.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1269,190.5,1269</points>
<connection>
<GID>164</GID>
<name>IN_B_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1270.5,189.5,1270.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1268,189.5,1268.5</points>
<intersection>1268 1</intersection>
<intersection>1268.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1268,190.5,1268</points>
<connection>
<GID>164</GID>
<name>IN_B_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1268.5,189.5,1268.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1266.5,189.5,1267</points>
<intersection>1266.5 2</intersection>
<intersection>1267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1267,190.5,1267</points>
<connection>
<GID>164</GID>
<name>IN_B_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1266.5,189.5,1266.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1264.5,189.5,1266</points>
<intersection>1264.5 2</intersection>
<intersection>1266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1266,190.5,1266</points>
<connection>
<GID>164</GID>
<name>IN_B_3</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1264.5,189.5,1264.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1262,189.5,1262.5</points>
<intersection>1262 1</intersection>
<intersection>1262.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1262,190.5,1262</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1262.5,189.5,1262.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1260.5,189.5,1261</points>
<intersection>1260.5 2</intersection>
<intersection>1261 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1261,190.5,1261</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1260.5,189.5,1260.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,1258.5,189.5,1260</points>
<intersection>1258.5 2</intersection>
<intersection>1260 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189.5,1260,190.5,1260</points>
<connection>
<GID>164</GID>
<name>IN_2</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1258.5,189.5,1258.5</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,1256.5,190,1259</points>
<intersection>1256.5 2</intersection>
<intersection>1259 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,1259,190.5,1259</points>
<connection>
<GID>164</GID>
<name>IN_3</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>188.5,1256.5,190,1256.5</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1299,262,1299</points>
<connection>
<GID>761</GID>
<name>IN_15</name></connection>
<connection>
<GID>763</GID>
<name>OUT_15</name></connection>
<intersection>258 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,1266,258,1299</points>
<connection>
<GID>762</GID>
<name>OUT_0</name></connection>
<intersection>1299 1</intersection></vsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1298,262,1298</points>
<connection>
<GID>761</GID>
<name>IN_14</name></connection>
<connection>
<GID>763</GID>
<name>OUT_14</name></connection>
<intersection>258 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,1267,258,1298</points>
<connection>
<GID>762</GID>
<name>OUT_1</name></connection>
<intersection>1298 1</intersection></vsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1297,262,1297</points>
<connection>
<GID>761</GID>
<name>IN_13</name></connection>
<connection>
<GID>763</GID>
<name>OUT_13</name></connection>
<intersection>258 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>258,1268,258,1297</points>
<connection>
<GID>762</GID>
<name>OUT_2</name></connection>
<intersection>1297 1</intersection></vsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1296,262,1296</points>
<connection>
<GID>761</GID>
<name>IN_12</name></connection>
<connection>
<GID>763</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1295,262,1295</points>
<connection>
<GID>761</GID>
<name>IN_11</name></connection>
<connection>
<GID>763</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1294,262,1294</points>
<connection>
<GID>761</GID>
<name>IN_10</name></connection>
<connection>
<GID>763</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1293,262,1293</points>
<connection>
<GID>761</GID>
<name>IN_9</name></connection>
<connection>
<GID>763</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1292,262,1292</points>
<connection>
<GID>761</GID>
<name>IN_8</name></connection>
<connection>
<GID>763</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1291,262,1291</points>
<connection>
<GID>761</GID>
<name>IN_7</name></connection>
<connection>
<GID>763</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1289,262,1289</points>
<connection>
<GID>761</GID>
<name>IN_5</name></connection>
<connection>
<GID>763</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1290,262,1290</points>
<connection>
<GID>761</GID>
<name>IN_6</name></connection>
<connection>
<GID>763</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>748</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1285,274.5,1285</points>
<connection>
<GID>761</GID>
<name>OUT_1</name></connection>
<connection>
<GID>296</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1288,262,1288</points>
<connection>
<GID>761</GID>
<name>IN_4</name></connection>
<connection>
<GID>763</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1286,262,1286</points>
<connection>
<GID>761</GID>
<name>IN_2</name></connection>
<connection>
<GID>763</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1287,262,1287</points>
<connection>
<GID>761</GID>
<name>IN_3</name></connection>
<connection>
<GID>763</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1285,262,1285</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<connection>
<GID>763</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258,1284,262,1284</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<connection>
<GID>763</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,1252,196.5,1256</points>
<connection>
<GID>164</GID>
<name>A_less_B</name></connection>
<intersection>1252 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,1252,254,1252</points>
<intersection>196.5 0</intersection>
<intersection>254 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>254,1252,254,1266</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>1252 1</intersection></vsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,1251,194.5,1256</points>
<connection>
<GID>164</GID>
<name>A_equal_B</name></connection>
<intersection>1251 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,1251,253,1251</points>
<intersection>194.5 0</intersection>
<intersection>253 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>253,1251,253,1267</points>
<intersection>1251 1</intersection>
<intersection>1267 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>253,1267,254,1267</points>
<connection>
<GID>762</GID>
<name>IN_1</name></connection>
<intersection>253 2</intersection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192.5,1250,192.5,1256</points>
<connection>
<GID>164</GID>
<name>A_greater_B</name></connection>
<intersection>1250 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192.5,1250,252,1250</points>
<intersection>192.5 0</intersection>
<intersection>252 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>252,1250,252,1268</points>
<intersection>1250 1</intersection>
<intersection>1268 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>252,1268,254,1268</points>
<connection>
<GID>762</GID>
<name>IN_2</name></connection>
<intersection>252 2</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,1300.5,264,1307</points>
<connection>
<GID>761</GID>
<name>ENABLE_0</name></connection>
<intersection>1307 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>256,1307,264,1307</points>
<connection>
<GID>702</GID>
<name>N_in1</name></connection>
<intersection>256 10</intersection>
<intersection>264 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>256,1307,256,1314</points>
<intersection>1307 9</intersection>
<intersection>1314 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>256,1314,261.5,1314</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>256 10</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253,1282,253,1307</points>
<intersection>1282 4</intersection>
<intersection>1300.5 5</intersection>
<intersection>1307 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>253,1282,256,1282</points>
<intersection>253 0</intersection>
<intersection>256 6</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>253,1300.5,256,1300.5</points>
<connection>
<GID>763</GID>
<name>ENABLE_0</name></connection>
<intersection>253 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>256,1278.5,256,1282</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>1282 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>253,1307,255,1307</points>
<connection>
<GID>702</GID>
<name>N_in0</name></connection>
<intersection>253 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,1270.5,256,1274.5</points>
<connection>
<GID>762</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1293,274.5,1293</points>
<connection>
<GID>761</GID>
<name>OUT_9</name></connection>
<connection>
<GID>272</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1292,268,1292</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1291,274.5,1291</points>
<connection>
<GID>761</GID>
<name>OUT_7</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1290,268,1290</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>761</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,1289,274.5,1289</points>
<connection>
<GID>761</GID>
<name>OUT_5</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-382.81,3701.51,1171.19,2686.51</PageViewport></page 2>
<page 3>
<PageViewport>-343.354,4254.68,1210.65,3239.68</PageViewport></page 3>
<page 4>
<PageViewport>-124.938,1792.26,1429.06,777.261</PageViewport></page 4>
<page 5>
<PageViewport>-296.679,2066.05,1257.32,1051.05</PageViewport></page 5>
<page 6>
<PageViewport>-251.668,4069.93,1302.33,3054.93</PageViewport></page 6>
<page 7>
<PageViewport>-251.668,4069.93,1302.33,3054.93</PageViewport></page 7>
<page 8>
<PageViewport>-251.668,4069.93,1302.33,3054.93</PageViewport></page 8>
<page 9>
<PageViewport>-251.668,4069.93,1302.33,3054.93</PageViewport></page 9></circuit>